module dadda_tree(
    input logic[31:0] opA,
    input logic[31:0] opB,
    output logic[63:0] row_top,
    output logic[63:0] row_bot
);

logic [31:0] comb[32];

genvar i, j;
for(i = 0; i < 32; ++i) begin
    for(j = 0; j < 32; ++j) begin
        assign comb[i][j] = opB[i] & opA[j];
    end
end
// stage 8 begin ======================================================================================================= 
logic S_s8_28_0, C_s8_28_0;
HA HA_s8_280(.A_i(comb[0][28]), .B_i(comb[1][27]), .S_o(S_s8_28_0), .c_out(C_s8_28_0));
logic S_s8_29_0, C_s8_29_0;
FA FA_s8_29_0(.A_i(comb[0][29]), .B_i(comb[1][28]), .c_in(comb[2][27]), .S_o(S_s8_29_0), .c_out(C_s8_29_0));
logic S_s8_29_1, C_s8_29_1;
HA HA_s8_291(.A_i(comb[3][26]), .B_i(comb[4][25]), .S_o(S_s8_29_1), .c_out(C_s8_29_1));
logic S_s8_30_0, C_s8_30_0;
FA FA_s8_30_0(.A_i(comb[0][30]), .B_i(comb[1][29]), .c_in(comb[2][28]), .S_o(S_s8_30_0), .c_out(C_s8_30_0));
logic S_s8_30_1, C_s8_30_1;
FA FA_s8_30_1(.A_i(comb[3][27]), .B_i(comb[4][26]), .c_in(comb[5][25]), .S_o(S_s8_30_1), .c_out(C_s8_30_1));
logic S_s8_30_2, C_s8_30_2;
HA HA_s8_302(.A_i(comb[6][24]), .B_i(comb[7][23]), .S_o(S_s8_30_2), .c_out(C_s8_30_2));
logic S_s8_31_0, C_s8_31_0;
FA FA_s8_31_0(.A_i(comb[0][31]), .B_i(comb[1][30]), .c_in(comb[2][29]), .S_o(S_s8_31_0), .c_out(C_s8_31_0));
logic S_s8_31_1, C_s8_31_1;
FA FA_s8_31_1(.A_i(comb[3][28]), .B_i(comb[4][27]), .c_in(comb[5][26]), .S_o(S_s8_31_1), .c_out(C_s8_31_1));
logic S_s8_31_2, C_s8_31_2;
FA FA_s8_31_2(.A_i(comb[6][25]), .B_i(comb[7][24]), .c_in(comb[8][23]), .S_o(S_s8_31_2), .c_out(C_s8_31_2));
logic S_s8_31_3, C_s8_31_3;
HA HA_s8_313(.A_i(comb[9][22]), .B_i(comb[10][21]), .S_o(S_s8_31_3), .c_out(C_s8_31_3));
logic S_s8_32_0, C_s8_32_0;
FA FA_s8_32_0(.A_i(comb[1][31]), .B_i(comb[2][30]), .c_in(comb[3][29]), .S_o(S_s8_32_0), .c_out(C_s8_32_0));
logic S_s8_32_1, C_s8_32_1;
FA FA_s8_32_1(.A_i(comb[4][28]), .B_i(comb[5][27]), .c_in(comb[6][26]), .S_o(S_s8_32_1), .c_out(C_s8_32_1));
logic S_s8_32_2, C_s8_32_2;
FA FA_s8_32_2(.A_i(comb[7][25]), .B_i(comb[8][24]), .c_in(comb[9][23]), .S_o(S_s8_32_2), .c_out(C_s8_32_2));
logic S_s8_32_3, C_s8_32_3;
HA HA_s8_323(.A_i(comb[10][22]), .B_i(comb[11][21]), .S_o(S_s8_32_3), .c_out(C_s8_32_3));
logic S_s8_33_0, C_s8_33_0;
FA FA_s8_33_0(.A_i(comb[2][31]), .B_i(comb[3][30]), .c_in(comb[4][29]), .S_o(S_s8_33_0), .c_out(C_s8_33_0));
logic S_s8_33_1, C_s8_33_1;
FA FA_s8_33_1(.A_i(comb[5][28]), .B_i(comb[6][27]), .c_in(comb[7][26]), .S_o(S_s8_33_1), .c_out(C_s8_33_1));
logic S_s8_33_2, C_s8_33_2;
FA FA_s8_33_2(.A_i(comb[8][25]), .B_i(comb[9][24]), .c_in(comb[10][23]), .S_o(S_s8_33_2), .c_out(C_s8_33_2));
logic S_s8_34_0, C_s8_34_0;
FA FA_s8_34_0(.A_i(comb[3][31]), .B_i(comb[4][30]), .c_in(comb[5][29]), .S_o(S_s8_34_0), .c_out(C_s8_34_0));
logic S_s8_34_1, C_s8_34_1;
FA FA_s8_34_1(.A_i(comb[6][28]), .B_i(comb[7][27]), .c_in(comb[8][26]), .S_o(S_s8_34_1), .c_out(C_s8_34_1));
logic S_s8_35_0, C_s8_35_0;
FA FA_s8_35_0(.A_i(comb[4][31]), .B_i(comb[5][30]), .c_in(comb[6][29]), .S_o(S_s8_35_0), .c_out(C_s8_35_0));
// stage 8 end ======================================================================================================= 

// stage 7 begin ======================================================================================================= 
logic S_s7_19_0, C_s7_19_0;
HA HA_s7_190(.A_i(comb[0][19]), .B_i(comb[1][18]), .S_o(S_s7_19_0), .c_out(C_s7_19_0));
logic S_s7_20_0, C_s7_20_0;
FA FA_s7_20_0(.A_i(comb[0][20]), .B_i(comb[1][19]), .c_in(comb[2][18]), .S_o(S_s7_20_0), .c_out(C_s7_20_0));
logic S_s7_20_1, C_s7_20_1;
HA HA_s7_201(.A_i(comb[3][17]), .B_i(comb[4][16]), .S_o(S_s7_20_1), .c_out(C_s7_20_1));
logic S_s7_21_0, C_s7_21_0;
FA FA_s7_21_0(.A_i(comb[0][21]), .B_i(comb[1][20]), .c_in(comb[2][19]), .S_o(S_s7_21_0), .c_out(C_s7_21_0));
logic S_s7_21_1, C_s7_21_1;
FA FA_s7_21_1(.A_i(comb[3][18]), .B_i(comb[4][17]), .c_in(comb[5][16]), .S_o(S_s7_21_1), .c_out(C_s7_21_1));
logic S_s7_21_2, C_s7_21_2;
HA HA_s7_212(.A_i(comb[6][15]), .B_i(comb[7][14]), .S_o(S_s7_21_2), .c_out(C_s7_21_2));
logic S_s7_22_0, C_s7_22_0;
FA FA_s7_22_0(.A_i(comb[0][22]), .B_i(comb[1][21]), .c_in(comb[2][20]), .S_o(S_s7_22_0), .c_out(C_s7_22_0));
logic S_s7_22_1, C_s7_22_1;
FA FA_s7_22_1(.A_i(comb[3][19]), .B_i(comb[4][18]), .c_in(comb[5][17]), .S_o(S_s7_22_1), .c_out(C_s7_22_1));
logic S_s7_22_2, C_s7_22_2;
FA FA_s7_22_2(.A_i(comb[6][16]), .B_i(comb[7][15]), .c_in(comb[8][14]), .S_o(S_s7_22_2), .c_out(C_s7_22_2));
logic S_s7_22_3, C_s7_22_3;
HA HA_s7_223(.A_i(comb[9][13]), .B_i(comb[10][12]), .S_o(S_s7_22_3), .c_out(C_s7_22_3));
logic S_s7_23_0, C_s7_23_0;
FA FA_s7_23_0(.A_i(comb[0][23]), .B_i(comb[1][22]), .c_in(comb[2][21]), .S_o(S_s7_23_0), .c_out(C_s7_23_0));
logic S_s7_23_1, C_s7_23_1;
FA FA_s7_23_1(.A_i(comb[3][20]), .B_i(comb[4][19]), .c_in(comb[5][18]), .S_o(S_s7_23_1), .c_out(C_s7_23_1));
logic S_s7_23_2, C_s7_23_2;
FA FA_s7_23_2(.A_i(comb[6][17]), .B_i(comb[7][16]), .c_in(comb[8][15]), .S_o(S_s7_23_2), .c_out(C_s7_23_2));
logic S_s7_23_3, C_s7_23_3;
FA FA_s7_23_3(.A_i(comb[9][14]), .B_i(comb[10][13]), .c_in(comb[11][12]), .S_o(S_s7_23_3), .c_out(C_s7_23_3));
logic S_s7_23_4, C_s7_23_4;
HA HA_s7_234(.A_i(comb[12][11]), .B_i(comb[13][10]), .S_o(S_s7_23_4), .c_out(C_s7_23_4));
logic S_s7_24_0, C_s7_24_0;
FA FA_s7_24_0(.A_i(comb[0][24]), .B_i(comb[1][23]), .c_in(comb[2][22]), .S_o(S_s7_24_0), .c_out(C_s7_24_0));
logic S_s7_24_1, C_s7_24_1;
FA FA_s7_24_1(.A_i(comb[3][21]), .B_i(comb[4][20]), .c_in(comb[5][19]), .S_o(S_s7_24_1), .c_out(C_s7_24_1));
logic S_s7_24_2, C_s7_24_2;
FA FA_s7_24_2(.A_i(comb[6][18]), .B_i(comb[7][17]), .c_in(comb[8][16]), .S_o(S_s7_24_2), .c_out(C_s7_24_2));
logic S_s7_24_3, C_s7_24_3;
FA FA_s7_24_3(.A_i(comb[9][15]), .B_i(comb[10][14]), .c_in(comb[11][13]), .S_o(S_s7_24_3), .c_out(C_s7_24_3));
logic S_s7_24_4, C_s7_24_4;
FA FA_s7_24_4(.A_i(comb[12][12]), .B_i(comb[13][11]), .c_in(comb[14][10]), .S_o(S_s7_24_4), .c_out(C_s7_24_4));
logic S_s7_24_5, C_s7_24_5;
HA HA_s7_245(.A_i(comb[15][9]), .B_i(comb[16][8]), .S_o(S_s7_24_5), .c_out(C_s7_24_5));
logic S_s7_25_0, C_s7_25_0;
FA FA_s7_25_0(.A_i(comb[0][25]), .B_i(comb[1][24]), .c_in(comb[2][23]), .S_o(S_s7_25_0), .c_out(C_s7_25_0));
logic S_s7_25_1, C_s7_25_1;
FA FA_s7_25_1(.A_i(comb[3][22]), .B_i(comb[4][21]), .c_in(comb[5][20]), .S_o(S_s7_25_1), .c_out(C_s7_25_1));
logic S_s7_25_2, C_s7_25_2;
FA FA_s7_25_2(.A_i(comb[6][19]), .B_i(comb[7][18]), .c_in(comb[8][17]), .S_o(S_s7_25_2), .c_out(C_s7_25_2));
logic S_s7_25_3, C_s7_25_3;
FA FA_s7_25_3(.A_i(comb[9][16]), .B_i(comb[10][15]), .c_in(comb[11][14]), .S_o(S_s7_25_3), .c_out(C_s7_25_3));
logic S_s7_25_4, C_s7_25_4;
FA FA_s7_25_4(.A_i(comb[12][13]), .B_i(comb[13][12]), .c_in(comb[14][11]), .S_o(S_s7_25_4), .c_out(C_s7_25_4));
logic S_s7_25_5, C_s7_25_5;
FA FA_s7_25_5(.A_i(comb[15][10]), .B_i(comb[16][9]), .c_in(comb[17][8]), .S_o(S_s7_25_5), .c_out(C_s7_25_5));
logic S_s7_25_6, C_s7_25_6;
HA HA_s7_256(.A_i(comb[18][7]), .B_i(comb[19][6]), .S_o(S_s7_25_6), .c_out(C_s7_25_6));
logic S_s7_26_0, C_s7_26_0;
FA FA_s7_26_0(.A_i(comb[0][26]), .B_i(comb[1][25]), .c_in(comb[2][24]), .S_o(S_s7_26_0), .c_out(C_s7_26_0));
logic S_s7_26_1, C_s7_26_1;
FA FA_s7_26_1(.A_i(comb[3][23]), .B_i(comb[4][22]), .c_in(comb[5][21]), .S_o(S_s7_26_1), .c_out(C_s7_26_1));
logic S_s7_26_2, C_s7_26_2;
FA FA_s7_26_2(.A_i(comb[6][20]), .B_i(comb[7][19]), .c_in(comb[8][18]), .S_o(S_s7_26_2), .c_out(C_s7_26_2));
logic S_s7_26_3, C_s7_26_3;
FA FA_s7_26_3(.A_i(comb[9][17]), .B_i(comb[10][16]), .c_in(comb[11][15]), .S_o(S_s7_26_3), .c_out(C_s7_26_3));
logic S_s7_26_4, C_s7_26_4;
FA FA_s7_26_4(.A_i(comb[12][14]), .B_i(comb[13][13]), .c_in(comb[14][12]), .S_o(S_s7_26_4), .c_out(C_s7_26_4));
logic S_s7_26_5, C_s7_26_5;
FA FA_s7_26_5(.A_i(comb[15][11]), .B_i(comb[16][10]), .c_in(comb[17][9]), .S_o(S_s7_26_5), .c_out(C_s7_26_5));
logic S_s7_26_6, C_s7_26_6;
FA FA_s7_26_6(.A_i(comb[18][8]), .B_i(comb[19][7]), .c_in(comb[20][6]), .S_o(S_s7_26_6), .c_out(C_s7_26_6));
logic S_s7_26_7, C_s7_26_7;
HA HA_s7_267(.A_i(comb[21][5]), .B_i(comb[22][4]), .S_o(S_s7_26_7), .c_out(C_s7_26_7));
logic S_s7_27_0, C_s7_27_0;
FA FA_s7_27_0(.A_i(comb[0][27]), .B_i(comb[1][26]), .c_in(comb[2][25]), .S_o(S_s7_27_0), .c_out(C_s7_27_0));
logic S_s7_27_1, C_s7_27_1;
FA FA_s7_27_1(.A_i(comb[3][24]), .B_i(comb[4][23]), .c_in(comb[5][22]), .S_o(S_s7_27_1), .c_out(C_s7_27_1));
logic S_s7_27_2, C_s7_27_2;
FA FA_s7_27_2(.A_i(comb[6][21]), .B_i(comb[7][20]), .c_in(comb[8][19]), .S_o(S_s7_27_2), .c_out(C_s7_27_2));
logic S_s7_27_3, C_s7_27_3;
FA FA_s7_27_3(.A_i(comb[9][18]), .B_i(comb[10][17]), .c_in(comb[11][16]), .S_o(S_s7_27_3), .c_out(C_s7_27_3));
logic S_s7_27_4, C_s7_27_4;
FA FA_s7_27_4(.A_i(comb[12][15]), .B_i(comb[13][14]), .c_in(comb[14][13]), .S_o(S_s7_27_4), .c_out(C_s7_27_4));
logic S_s7_27_5, C_s7_27_5;
FA FA_s7_27_5(.A_i(comb[15][12]), .B_i(comb[16][11]), .c_in(comb[17][10]), .S_o(S_s7_27_5), .c_out(C_s7_27_5));
logic S_s7_27_6, C_s7_27_6;
FA FA_s7_27_6(.A_i(comb[18][9]), .B_i(comb[19][8]), .c_in(comb[20][7]), .S_o(S_s7_27_6), .c_out(C_s7_27_6));
logic S_s7_27_7, C_s7_27_7;
FA FA_s7_27_7(.A_i(comb[21][6]), .B_i(comb[22][5]), .c_in(comb[23][4]), .S_o(S_s7_27_7), .c_out(C_s7_27_7));
logic S_s7_27_8, C_s7_27_8;
HA HA_s7_278(.A_i(comb[24][3]), .B_i(comb[25][2]), .S_o(S_s7_27_8), .c_out(C_s7_27_8));
logic S_s7_28_0, C_s7_28_0;
FA FA_s7_28_0(.A_i(S_s8_28_0), .B_i(comb[2][26]), .c_in(comb[3][25]), .S_o(S_s7_28_0), .c_out(C_s7_28_0));
logic S_s7_28_1, C_s7_28_1;
FA FA_s7_28_1(.A_i(comb[4][24]), .B_i(comb[5][23]), .c_in(comb[6][22]), .S_o(S_s7_28_1), .c_out(C_s7_28_1));
logic S_s7_28_2, C_s7_28_2;
FA FA_s7_28_2(.A_i(comb[7][21]), .B_i(comb[8][20]), .c_in(comb[9][19]), .S_o(S_s7_28_2), .c_out(C_s7_28_2));
logic S_s7_28_3, C_s7_28_3;
FA FA_s7_28_3(.A_i(comb[10][18]), .B_i(comb[11][17]), .c_in(comb[12][16]), .S_o(S_s7_28_3), .c_out(C_s7_28_3));
logic S_s7_28_4, C_s7_28_4;
FA FA_s7_28_4(.A_i(comb[13][15]), .B_i(comb[14][14]), .c_in(comb[15][13]), .S_o(S_s7_28_4), .c_out(C_s7_28_4));
logic S_s7_28_5, C_s7_28_5;
FA FA_s7_28_5(.A_i(comb[16][12]), .B_i(comb[17][11]), .c_in(comb[18][10]), .S_o(S_s7_28_5), .c_out(C_s7_28_5));
logic S_s7_28_6, C_s7_28_6;
FA FA_s7_28_6(.A_i(comb[19][9]), .B_i(comb[20][8]), .c_in(comb[21][7]), .S_o(S_s7_28_6), .c_out(C_s7_28_6));
logic S_s7_28_7, C_s7_28_7;
FA FA_s7_28_7(.A_i(comb[22][6]), .B_i(comb[23][5]), .c_in(comb[24][4]), .S_o(S_s7_28_7), .c_out(C_s7_28_7));
logic S_s7_28_8, C_s7_28_8;
FA FA_s7_28_8(.A_i(comb[25][3]), .B_i(comb[26][2]), .c_in(comb[27][1]), .S_o(S_s7_28_8), .c_out(C_s7_28_8));
logic S_s7_29_0, C_s7_29_0;
FA FA_s7_29_0(.A_i(S_s8_29_1), .B_i(S_s8_29_0), .c_in(C_s8_28_0), .S_o(S_s7_29_0), .c_out(C_s7_29_0));
logic S_s7_29_1, C_s7_29_1;
FA FA_s7_29_1(.A_i(comb[5][24]), .B_i(comb[6][23]), .c_in(comb[7][22]), .S_o(S_s7_29_1), .c_out(C_s7_29_1));
logic S_s7_29_2, C_s7_29_2;
FA FA_s7_29_2(.A_i(comb[8][21]), .B_i(comb[9][20]), .c_in(comb[10][19]), .S_o(S_s7_29_2), .c_out(C_s7_29_2));
logic S_s7_29_3, C_s7_29_3;
FA FA_s7_29_3(.A_i(comb[11][18]), .B_i(comb[12][17]), .c_in(comb[13][16]), .S_o(S_s7_29_3), .c_out(C_s7_29_3));
logic S_s7_29_4, C_s7_29_4;
FA FA_s7_29_4(.A_i(comb[14][15]), .B_i(comb[15][14]), .c_in(comb[16][13]), .S_o(S_s7_29_4), .c_out(C_s7_29_4));
logic S_s7_29_5, C_s7_29_5;
FA FA_s7_29_5(.A_i(comb[17][12]), .B_i(comb[18][11]), .c_in(comb[19][10]), .S_o(S_s7_29_5), .c_out(C_s7_29_5));
logic S_s7_29_6, C_s7_29_6;
FA FA_s7_29_6(.A_i(comb[20][9]), .B_i(comb[21][8]), .c_in(comb[22][7]), .S_o(S_s7_29_6), .c_out(C_s7_29_6));
logic S_s7_29_7, C_s7_29_7;
FA FA_s7_29_7(.A_i(comb[23][6]), .B_i(comb[24][5]), .c_in(comb[25][4]), .S_o(S_s7_29_7), .c_out(C_s7_29_7));
logic S_s7_29_8, C_s7_29_8;
FA FA_s7_29_8(.A_i(comb[26][3]), .B_i(comb[27][2]), .c_in(comb[28][1]), .S_o(S_s7_29_8), .c_out(C_s7_29_8));
logic S_s7_30_0, C_s7_30_0;
FA FA_s7_30_0(.A_i(S_s8_30_2), .B_i(S_s8_30_1), .c_in(S_s8_30_0), .S_o(S_s7_30_0), .c_out(C_s7_30_0));
logic S_s7_30_1, C_s7_30_1;
FA FA_s7_30_1(.A_i(C_s8_29_1), .B_i(C_s8_29_0), .c_in(comb[8][22]), .S_o(S_s7_30_1), .c_out(C_s7_30_1));
logic S_s7_30_2, C_s7_30_2;
FA FA_s7_30_2(.A_i(comb[9][21]), .B_i(comb[10][20]), .c_in(comb[11][19]), .S_o(S_s7_30_2), .c_out(C_s7_30_2));
logic S_s7_30_3, C_s7_30_3;
FA FA_s7_30_3(.A_i(comb[12][18]), .B_i(comb[13][17]), .c_in(comb[14][16]), .S_o(S_s7_30_3), .c_out(C_s7_30_3));
logic S_s7_30_4, C_s7_30_4;
FA FA_s7_30_4(.A_i(comb[15][15]), .B_i(comb[16][14]), .c_in(comb[17][13]), .S_o(S_s7_30_4), .c_out(C_s7_30_4));
logic S_s7_30_5, C_s7_30_5;
FA FA_s7_30_5(.A_i(comb[18][12]), .B_i(comb[19][11]), .c_in(comb[20][10]), .S_o(S_s7_30_5), .c_out(C_s7_30_5));
logic S_s7_30_6, C_s7_30_6;
FA FA_s7_30_6(.A_i(comb[21][9]), .B_i(comb[22][8]), .c_in(comb[23][7]), .S_o(S_s7_30_6), .c_out(C_s7_30_6));
logic S_s7_30_7, C_s7_30_7;
FA FA_s7_30_7(.A_i(comb[24][6]), .B_i(comb[25][5]), .c_in(comb[26][4]), .S_o(S_s7_30_7), .c_out(C_s7_30_7));
logic S_s7_30_8, C_s7_30_8;
FA FA_s7_30_8(.A_i(comb[27][3]), .B_i(comb[28][2]), .c_in(comb[29][1]), .S_o(S_s7_30_8), .c_out(C_s7_30_8));
logic S_s7_31_0, C_s7_31_0;
FA FA_s7_31_0(.A_i(S_s8_31_3), .B_i(S_s8_31_2), .c_in(S_s8_31_1), .S_o(S_s7_31_0), .c_out(C_s7_31_0));
logic S_s7_31_1, C_s7_31_1;
FA FA_s7_31_1(.A_i(S_s8_31_0), .B_i(C_s8_30_2), .c_in(C_s8_30_1), .S_o(S_s7_31_1), .c_out(C_s7_31_1));
logic S_s7_31_2, C_s7_31_2;
FA FA_s7_31_2(.A_i(C_s8_30_0), .B_i(comb[11][20]), .c_in(comb[12][19]), .S_o(S_s7_31_2), .c_out(C_s7_31_2));
logic S_s7_31_3, C_s7_31_3;
FA FA_s7_31_3(.A_i(comb[13][18]), .B_i(comb[14][17]), .c_in(comb[15][16]), .S_o(S_s7_31_3), .c_out(C_s7_31_3));
logic S_s7_31_4, C_s7_31_4;
FA FA_s7_31_4(.A_i(comb[16][15]), .B_i(comb[17][14]), .c_in(comb[18][13]), .S_o(S_s7_31_4), .c_out(C_s7_31_4));
logic S_s7_31_5, C_s7_31_5;
FA FA_s7_31_5(.A_i(comb[19][12]), .B_i(comb[20][11]), .c_in(comb[21][10]), .S_o(S_s7_31_5), .c_out(C_s7_31_5));
logic S_s7_31_6, C_s7_31_6;
FA FA_s7_31_6(.A_i(comb[22][9]), .B_i(comb[23][8]), .c_in(comb[24][7]), .S_o(S_s7_31_6), .c_out(C_s7_31_6));
logic S_s7_31_7, C_s7_31_7;
FA FA_s7_31_7(.A_i(comb[25][6]), .B_i(comb[26][5]), .c_in(comb[27][4]), .S_o(S_s7_31_7), .c_out(C_s7_31_7));
logic S_s7_31_8, C_s7_31_8;
FA FA_s7_31_8(.A_i(comb[28][3]), .B_i(comb[29][2]), .c_in(comb[30][1]), .S_o(S_s7_31_8), .c_out(C_s7_31_8));
logic S_s7_32_0, C_s7_32_0;
FA FA_s7_32_0(.A_i(S_s8_32_3), .B_i(S_s8_32_2), .c_in(S_s8_32_1), .S_o(S_s7_32_0), .c_out(C_s7_32_0));
logic S_s7_32_1, C_s7_32_1;
FA FA_s7_32_1(.A_i(S_s8_32_0), .B_i(C_s8_31_3), .c_in(C_s8_31_2), .S_o(S_s7_32_1), .c_out(C_s7_32_1));
logic S_s7_32_2, C_s7_32_2;
FA FA_s7_32_2(.A_i(C_s8_31_1), .B_i(C_s8_31_0), .c_in(comb[12][20]), .S_o(S_s7_32_2), .c_out(C_s7_32_2));
logic S_s7_32_3, C_s7_32_3;
FA FA_s7_32_3(.A_i(comb[13][19]), .B_i(comb[14][18]), .c_in(comb[15][17]), .S_o(S_s7_32_3), .c_out(C_s7_32_3));
logic S_s7_32_4, C_s7_32_4;
FA FA_s7_32_4(.A_i(comb[16][16]), .B_i(comb[17][15]), .c_in(comb[18][14]), .S_o(S_s7_32_4), .c_out(C_s7_32_4));
logic S_s7_32_5, C_s7_32_5;
FA FA_s7_32_5(.A_i(comb[19][13]), .B_i(comb[20][12]), .c_in(comb[21][11]), .S_o(S_s7_32_5), .c_out(C_s7_32_5));
logic S_s7_32_6, C_s7_32_6;
FA FA_s7_32_6(.A_i(comb[22][10]), .B_i(comb[23][9]), .c_in(comb[24][8]), .S_o(S_s7_32_6), .c_out(C_s7_32_6));
logic S_s7_32_7, C_s7_32_7;
FA FA_s7_32_7(.A_i(comb[25][7]), .B_i(comb[26][6]), .c_in(comb[27][5]), .S_o(S_s7_32_7), .c_out(C_s7_32_7));
logic S_s7_32_8, C_s7_32_8;
FA FA_s7_32_8(.A_i(comb[28][4]), .B_i(comb[29][3]), .c_in(comb[30][2]), .S_o(S_s7_32_8), .c_out(C_s7_32_8));
logic S_s7_33_0, C_s7_33_0;
FA FA_s7_33_0(.A_i(S_s8_33_2), .B_i(S_s8_33_1), .c_in(S_s8_33_0), .S_o(S_s7_33_0), .c_out(C_s7_33_0));
logic S_s7_33_1, C_s7_33_1;
FA FA_s7_33_1(.A_i(C_s8_32_3), .B_i(C_s8_32_2), .c_in(C_s8_32_1), .S_o(S_s7_33_1), .c_out(C_s7_33_1));
logic S_s7_33_2, C_s7_33_2;
FA FA_s7_33_2(.A_i(C_s8_32_0), .B_i(comb[11][22]), .c_in(comb[12][21]), .S_o(S_s7_33_2), .c_out(C_s7_33_2));
logic S_s7_33_3, C_s7_33_3;
FA FA_s7_33_3(.A_i(comb[13][20]), .B_i(comb[14][19]), .c_in(comb[15][18]), .S_o(S_s7_33_3), .c_out(C_s7_33_3));
logic S_s7_33_4, C_s7_33_4;
FA FA_s7_33_4(.A_i(comb[16][17]), .B_i(comb[17][16]), .c_in(comb[18][15]), .S_o(S_s7_33_4), .c_out(C_s7_33_4));
logic S_s7_33_5, C_s7_33_5;
FA FA_s7_33_5(.A_i(comb[19][14]), .B_i(comb[20][13]), .c_in(comb[21][12]), .S_o(S_s7_33_5), .c_out(C_s7_33_5));
logic S_s7_33_6, C_s7_33_6;
FA FA_s7_33_6(.A_i(comb[22][11]), .B_i(comb[23][10]), .c_in(comb[24][9]), .S_o(S_s7_33_6), .c_out(C_s7_33_6));
logic S_s7_33_7, C_s7_33_7;
FA FA_s7_33_7(.A_i(comb[25][8]), .B_i(comb[26][7]), .c_in(comb[27][6]), .S_o(S_s7_33_7), .c_out(C_s7_33_7));
logic S_s7_33_8, C_s7_33_8;
FA FA_s7_33_8(.A_i(comb[28][5]), .B_i(comb[29][4]), .c_in(comb[30][3]), .S_o(S_s7_33_8), .c_out(C_s7_33_8));
logic S_s7_34_0, C_s7_34_0;
FA FA_s7_34_0(.A_i(S_s8_34_1), .B_i(S_s8_34_0), .c_in(C_s8_33_2), .S_o(S_s7_34_0), .c_out(C_s7_34_0));
logic S_s7_34_1, C_s7_34_1;
FA FA_s7_34_1(.A_i(C_s8_33_1), .B_i(C_s8_33_0), .c_in(comb[9][25]), .S_o(S_s7_34_1), .c_out(C_s7_34_1));
logic S_s7_34_2, C_s7_34_2;
FA FA_s7_34_2(.A_i(comb[10][24]), .B_i(comb[11][23]), .c_in(comb[12][22]), .S_o(S_s7_34_2), .c_out(C_s7_34_2));
logic S_s7_34_3, C_s7_34_3;
FA FA_s7_34_3(.A_i(comb[13][21]), .B_i(comb[14][20]), .c_in(comb[15][19]), .S_o(S_s7_34_3), .c_out(C_s7_34_3));
logic S_s7_34_4, C_s7_34_4;
FA FA_s7_34_4(.A_i(comb[16][18]), .B_i(comb[17][17]), .c_in(comb[18][16]), .S_o(S_s7_34_4), .c_out(C_s7_34_4));
logic S_s7_34_5, C_s7_34_5;
FA FA_s7_34_5(.A_i(comb[19][15]), .B_i(comb[20][14]), .c_in(comb[21][13]), .S_o(S_s7_34_5), .c_out(C_s7_34_5));
logic S_s7_34_6, C_s7_34_6;
FA FA_s7_34_6(.A_i(comb[22][12]), .B_i(comb[23][11]), .c_in(comb[24][10]), .S_o(S_s7_34_6), .c_out(C_s7_34_6));
logic S_s7_34_7, C_s7_34_7;
FA FA_s7_34_7(.A_i(comb[25][9]), .B_i(comb[26][8]), .c_in(comb[27][7]), .S_o(S_s7_34_7), .c_out(C_s7_34_7));
logic S_s7_34_8, C_s7_34_8;
FA FA_s7_34_8(.A_i(comb[28][6]), .B_i(comb[29][5]), .c_in(comb[30][4]), .S_o(S_s7_34_8), .c_out(C_s7_34_8));
logic S_s7_35_0, C_s7_35_0;
FA FA_s7_35_0(.A_i(S_s8_35_0), .B_i(C_s8_34_1), .c_in(C_s8_34_0), .S_o(S_s7_35_0), .c_out(C_s7_35_0));
logic S_s7_35_1, C_s7_35_1;
FA FA_s7_35_1(.A_i(comb[7][28]), .B_i(comb[8][27]), .c_in(comb[9][26]), .S_o(S_s7_35_1), .c_out(C_s7_35_1));
logic S_s7_35_2, C_s7_35_2;
FA FA_s7_35_2(.A_i(comb[10][25]), .B_i(comb[11][24]), .c_in(comb[12][23]), .S_o(S_s7_35_2), .c_out(C_s7_35_2));
logic S_s7_35_3, C_s7_35_3;
FA FA_s7_35_3(.A_i(comb[13][22]), .B_i(comb[14][21]), .c_in(comb[15][20]), .S_o(S_s7_35_3), .c_out(C_s7_35_3));
logic S_s7_35_4, C_s7_35_4;
FA FA_s7_35_4(.A_i(comb[16][19]), .B_i(comb[17][18]), .c_in(comb[18][17]), .S_o(S_s7_35_4), .c_out(C_s7_35_4));
logic S_s7_35_5, C_s7_35_5;
FA FA_s7_35_5(.A_i(comb[19][16]), .B_i(comb[20][15]), .c_in(comb[21][14]), .S_o(S_s7_35_5), .c_out(C_s7_35_5));
logic S_s7_35_6, C_s7_35_6;
FA FA_s7_35_6(.A_i(comb[22][13]), .B_i(comb[23][12]), .c_in(comb[24][11]), .S_o(S_s7_35_6), .c_out(C_s7_35_6));
logic S_s7_35_7, C_s7_35_7;
FA FA_s7_35_7(.A_i(comb[25][10]), .B_i(comb[26][9]), .c_in(comb[27][8]), .S_o(S_s7_35_7), .c_out(C_s7_35_7));
logic S_s7_35_8, C_s7_35_8;
FA FA_s7_35_8(.A_i(comb[28][7]), .B_i(comb[29][6]), .c_in(comb[30][5]), .S_o(S_s7_35_8), .c_out(C_s7_35_8));
logic S_s7_36_0, C_s7_36_0;
FA FA_s7_36_0(.A_i(C_s8_35_0), .B_i(comb[5][31]), .c_in(comb[6][30]), .S_o(S_s7_36_0), .c_out(C_s7_36_0));
logic S_s7_36_1, C_s7_36_1;
FA FA_s7_36_1(.A_i(comb[7][29]), .B_i(comb[8][28]), .c_in(comb[9][27]), .S_o(S_s7_36_1), .c_out(C_s7_36_1));
logic S_s7_36_2, C_s7_36_2;
FA FA_s7_36_2(.A_i(comb[10][26]), .B_i(comb[11][25]), .c_in(comb[12][24]), .S_o(S_s7_36_2), .c_out(C_s7_36_2));
logic S_s7_36_3, C_s7_36_3;
FA FA_s7_36_3(.A_i(comb[13][23]), .B_i(comb[14][22]), .c_in(comb[15][21]), .S_o(S_s7_36_3), .c_out(C_s7_36_3));
logic S_s7_36_4, C_s7_36_4;
FA FA_s7_36_4(.A_i(comb[16][20]), .B_i(comb[17][19]), .c_in(comb[18][18]), .S_o(S_s7_36_4), .c_out(C_s7_36_4));
logic S_s7_36_5, C_s7_36_5;
FA FA_s7_36_5(.A_i(comb[19][17]), .B_i(comb[20][16]), .c_in(comb[21][15]), .S_o(S_s7_36_5), .c_out(C_s7_36_5));
logic S_s7_36_6, C_s7_36_6;
FA FA_s7_36_6(.A_i(comb[22][14]), .B_i(comb[23][13]), .c_in(comb[24][12]), .S_o(S_s7_36_6), .c_out(C_s7_36_6));
logic S_s7_36_7, C_s7_36_7;
FA FA_s7_36_7(.A_i(comb[25][11]), .B_i(comb[26][10]), .c_in(comb[27][9]), .S_o(S_s7_36_7), .c_out(C_s7_36_7));
logic S_s7_36_8, C_s7_36_8;
FA FA_s7_36_8(.A_i(comb[28][8]), .B_i(comb[29][7]), .c_in(comb[30][6]), .S_o(S_s7_36_8), .c_out(C_s7_36_8));
logic S_s7_37_0, C_s7_37_0;
FA FA_s7_37_0(.A_i(comb[6][31]), .B_i(comb[7][30]), .c_in(comb[8][29]), .S_o(S_s7_37_0), .c_out(C_s7_37_0));
logic S_s7_37_1, C_s7_37_1;
FA FA_s7_37_1(.A_i(comb[9][28]), .B_i(comb[10][27]), .c_in(comb[11][26]), .S_o(S_s7_37_1), .c_out(C_s7_37_1));
logic S_s7_37_2, C_s7_37_2;
FA FA_s7_37_2(.A_i(comb[12][25]), .B_i(comb[13][24]), .c_in(comb[14][23]), .S_o(S_s7_37_2), .c_out(C_s7_37_2));
logic S_s7_37_3, C_s7_37_3;
FA FA_s7_37_3(.A_i(comb[15][22]), .B_i(comb[16][21]), .c_in(comb[17][20]), .S_o(S_s7_37_3), .c_out(C_s7_37_3));
logic S_s7_37_4, C_s7_37_4;
FA FA_s7_37_4(.A_i(comb[18][19]), .B_i(comb[19][18]), .c_in(comb[20][17]), .S_o(S_s7_37_4), .c_out(C_s7_37_4));
logic S_s7_37_5, C_s7_37_5;
FA FA_s7_37_5(.A_i(comb[21][16]), .B_i(comb[22][15]), .c_in(comb[23][14]), .S_o(S_s7_37_5), .c_out(C_s7_37_5));
logic S_s7_37_6, C_s7_37_6;
FA FA_s7_37_6(.A_i(comb[24][13]), .B_i(comb[25][12]), .c_in(comb[26][11]), .S_o(S_s7_37_6), .c_out(C_s7_37_6));
logic S_s7_37_7, C_s7_37_7;
FA FA_s7_37_7(.A_i(comb[27][10]), .B_i(comb[28][9]), .c_in(comb[29][8]), .S_o(S_s7_37_7), .c_out(C_s7_37_7));
logic S_s7_38_0, C_s7_38_0;
FA FA_s7_38_0(.A_i(comb[7][31]), .B_i(comb[8][30]), .c_in(comb[9][29]), .S_o(S_s7_38_0), .c_out(C_s7_38_0));
logic S_s7_38_1, C_s7_38_1;
FA FA_s7_38_1(.A_i(comb[10][28]), .B_i(comb[11][27]), .c_in(comb[12][26]), .S_o(S_s7_38_1), .c_out(C_s7_38_1));
logic S_s7_38_2, C_s7_38_2;
FA FA_s7_38_2(.A_i(comb[13][25]), .B_i(comb[14][24]), .c_in(comb[15][23]), .S_o(S_s7_38_2), .c_out(C_s7_38_2));
logic S_s7_38_3, C_s7_38_3;
FA FA_s7_38_3(.A_i(comb[16][22]), .B_i(comb[17][21]), .c_in(comb[18][20]), .S_o(S_s7_38_3), .c_out(C_s7_38_3));
logic S_s7_38_4, C_s7_38_4;
FA FA_s7_38_4(.A_i(comb[19][19]), .B_i(comb[20][18]), .c_in(comb[21][17]), .S_o(S_s7_38_4), .c_out(C_s7_38_4));
logic S_s7_38_5, C_s7_38_5;
FA FA_s7_38_5(.A_i(comb[22][16]), .B_i(comb[23][15]), .c_in(comb[24][14]), .S_o(S_s7_38_5), .c_out(C_s7_38_5));
logic S_s7_38_6, C_s7_38_6;
FA FA_s7_38_6(.A_i(comb[25][13]), .B_i(comb[26][12]), .c_in(comb[27][11]), .S_o(S_s7_38_6), .c_out(C_s7_38_6));
logic S_s7_39_0, C_s7_39_0;
FA FA_s7_39_0(.A_i(comb[8][31]), .B_i(comb[9][30]), .c_in(comb[10][29]), .S_o(S_s7_39_0), .c_out(C_s7_39_0));
logic S_s7_39_1, C_s7_39_1;
FA FA_s7_39_1(.A_i(comb[11][28]), .B_i(comb[12][27]), .c_in(comb[13][26]), .S_o(S_s7_39_1), .c_out(C_s7_39_1));
logic S_s7_39_2, C_s7_39_2;
FA FA_s7_39_2(.A_i(comb[14][25]), .B_i(comb[15][24]), .c_in(comb[16][23]), .S_o(S_s7_39_2), .c_out(C_s7_39_2));
logic S_s7_39_3, C_s7_39_3;
FA FA_s7_39_3(.A_i(comb[17][22]), .B_i(comb[18][21]), .c_in(comb[19][20]), .S_o(S_s7_39_3), .c_out(C_s7_39_3));
logic S_s7_39_4, C_s7_39_4;
FA FA_s7_39_4(.A_i(comb[20][19]), .B_i(comb[21][18]), .c_in(comb[22][17]), .S_o(S_s7_39_4), .c_out(C_s7_39_4));
logic S_s7_39_5, C_s7_39_5;
FA FA_s7_39_5(.A_i(comb[23][16]), .B_i(comb[24][15]), .c_in(comb[25][14]), .S_o(S_s7_39_5), .c_out(C_s7_39_5));
logic S_s7_40_0, C_s7_40_0;
FA FA_s7_40_0(.A_i(comb[9][31]), .B_i(comb[10][30]), .c_in(comb[11][29]), .S_o(S_s7_40_0), .c_out(C_s7_40_0));
logic S_s7_40_1, C_s7_40_1;
FA FA_s7_40_1(.A_i(comb[12][28]), .B_i(comb[13][27]), .c_in(comb[14][26]), .S_o(S_s7_40_1), .c_out(C_s7_40_1));
logic S_s7_40_2, C_s7_40_2;
FA FA_s7_40_2(.A_i(comb[15][25]), .B_i(comb[16][24]), .c_in(comb[17][23]), .S_o(S_s7_40_2), .c_out(C_s7_40_2));
logic S_s7_40_3, C_s7_40_3;
FA FA_s7_40_3(.A_i(comb[18][22]), .B_i(comb[19][21]), .c_in(comb[20][20]), .S_o(S_s7_40_3), .c_out(C_s7_40_3));
logic S_s7_40_4, C_s7_40_4;
FA FA_s7_40_4(.A_i(comb[21][19]), .B_i(comb[22][18]), .c_in(comb[23][17]), .S_o(S_s7_40_4), .c_out(C_s7_40_4));
logic S_s7_41_0, C_s7_41_0;
FA FA_s7_41_0(.A_i(comb[10][31]), .B_i(comb[11][30]), .c_in(comb[12][29]), .S_o(S_s7_41_0), .c_out(C_s7_41_0));
logic S_s7_41_1, C_s7_41_1;
FA FA_s7_41_1(.A_i(comb[13][28]), .B_i(comb[14][27]), .c_in(comb[15][26]), .S_o(S_s7_41_1), .c_out(C_s7_41_1));
logic S_s7_41_2, C_s7_41_2;
FA FA_s7_41_2(.A_i(comb[16][25]), .B_i(comb[17][24]), .c_in(comb[18][23]), .S_o(S_s7_41_2), .c_out(C_s7_41_2));
logic S_s7_41_3, C_s7_41_3;
FA FA_s7_41_3(.A_i(comb[19][22]), .B_i(comb[20][21]), .c_in(comb[21][20]), .S_o(S_s7_41_3), .c_out(C_s7_41_3));
logic S_s7_42_0, C_s7_42_0;
FA FA_s7_42_0(.A_i(comb[11][31]), .B_i(comb[12][30]), .c_in(comb[13][29]), .S_o(S_s7_42_0), .c_out(C_s7_42_0));
logic S_s7_42_1, C_s7_42_1;
FA FA_s7_42_1(.A_i(comb[14][28]), .B_i(comb[15][27]), .c_in(comb[16][26]), .S_o(S_s7_42_1), .c_out(C_s7_42_1));
logic S_s7_42_2, C_s7_42_2;
FA FA_s7_42_2(.A_i(comb[17][25]), .B_i(comb[18][24]), .c_in(comb[19][23]), .S_o(S_s7_42_2), .c_out(C_s7_42_2));
logic S_s7_43_0, C_s7_43_0;
FA FA_s7_43_0(.A_i(comb[12][31]), .B_i(comb[13][30]), .c_in(comb[14][29]), .S_o(S_s7_43_0), .c_out(C_s7_43_0));
logic S_s7_43_1, C_s7_43_1;
FA FA_s7_43_1(.A_i(comb[15][28]), .B_i(comb[16][27]), .c_in(comb[17][26]), .S_o(S_s7_43_1), .c_out(C_s7_43_1));
logic S_s7_44_0, C_s7_44_0;
FA FA_s7_44_0(.A_i(comb[13][31]), .B_i(comb[14][30]), .c_in(comb[15][29]), .S_o(S_s7_44_0), .c_out(C_s7_44_0));
// stage 7 end ======================================================================================================= 

// stage 6 begin ======================================================================================================= 
logic S_s6_13_0, C_s6_13_0;
HA HA_s6_130(.A_i(comb[0][13]), .B_i(comb[1][12]), .S_o(S_s6_13_0), .c_out(C_s6_13_0));
logic S_s6_14_0, C_s6_14_0;
FA FA_s6_14_0(.A_i(comb[0][14]), .B_i(comb[1][13]), .c_in(comb[2][12]), .S_o(S_s6_14_0), .c_out(C_s6_14_0));
logic S_s6_14_1, C_s6_14_1;
HA HA_s6_141(.A_i(comb[3][11]), .B_i(comb[4][10]), .S_o(S_s6_14_1), .c_out(C_s6_14_1));
logic S_s6_15_0, C_s6_15_0;
FA FA_s6_15_0(.A_i(comb[0][15]), .B_i(comb[1][14]), .c_in(comb[2][13]), .S_o(S_s6_15_0), .c_out(C_s6_15_0));
logic S_s6_15_1, C_s6_15_1;
FA FA_s6_15_1(.A_i(comb[3][12]), .B_i(comb[4][11]), .c_in(comb[5][10]), .S_o(S_s6_15_1), .c_out(C_s6_15_1));
logic S_s6_15_2, C_s6_15_2;
HA HA_s6_152(.A_i(comb[6][9]), .B_i(comb[7][8]), .S_o(S_s6_15_2), .c_out(C_s6_15_2));
logic S_s6_16_0, C_s6_16_0;
FA FA_s6_16_0(.A_i(comb[0][16]), .B_i(comb[1][15]), .c_in(comb[2][14]), .S_o(S_s6_16_0), .c_out(C_s6_16_0));
logic S_s6_16_1, C_s6_16_1;
FA FA_s6_16_1(.A_i(comb[3][13]), .B_i(comb[4][12]), .c_in(comb[5][11]), .S_o(S_s6_16_1), .c_out(C_s6_16_1));
logic S_s6_16_2, C_s6_16_2;
FA FA_s6_16_2(.A_i(comb[6][10]), .B_i(comb[7][9]), .c_in(comb[8][8]), .S_o(S_s6_16_2), .c_out(C_s6_16_2));
logic S_s6_16_3, C_s6_16_3;
HA HA_s6_163(.A_i(comb[9][7]), .B_i(comb[10][6]), .S_o(S_s6_16_3), .c_out(C_s6_16_3));
logic S_s6_17_0, C_s6_17_0;
FA FA_s6_17_0(.A_i(comb[0][17]), .B_i(comb[1][16]), .c_in(comb[2][15]), .S_o(S_s6_17_0), .c_out(C_s6_17_0));
logic S_s6_17_1, C_s6_17_1;
FA FA_s6_17_1(.A_i(comb[3][14]), .B_i(comb[4][13]), .c_in(comb[5][12]), .S_o(S_s6_17_1), .c_out(C_s6_17_1));
logic S_s6_17_2, C_s6_17_2;
FA FA_s6_17_2(.A_i(comb[6][11]), .B_i(comb[7][10]), .c_in(comb[8][9]), .S_o(S_s6_17_2), .c_out(C_s6_17_2));
logic S_s6_17_3, C_s6_17_3;
FA FA_s6_17_3(.A_i(comb[9][8]), .B_i(comb[10][7]), .c_in(comb[11][6]), .S_o(S_s6_17_3), .c_out(C_s6_17_3));
logic S_s6_17_4, C_s6_17_4;
HA HA_s6_174(.A_i(comb[12][5]), .B_i(comb[13][4]), .S_o(S_s6_17_4), .c_out(C_s6_17_4));
logic S_s6_18_0, C_s6_18_0;
FA FA_s6_18_0(.A_i(comb[0][18]), .B_i(comb[1][17]), .c_in(comb[2][16]), .S_o(S_s6_18_0), .c_out(C_s6_18_0));
logic S_s6_18_1, C_s6_18_1;
FA FA_s6_18_1(.A_i(comb[3][15]), .B_i(comb[4][14]), .c_in(comb[5][13]), .S_o(S_s6_18_1), .c_out(C_s6_18_1));
logic S_s6_18_2, C_s6_18_2;
FA FA_s6_18_2(.A_i(comb[6][12]), .B_i(comb[7][11]), .c_in(comb[8][10]), .S_o(S_s6_18_2), .c_out(C_s6_18_2));
logic S_s6_18_3, C_s6_18_3;
FA FA_s6_18_3(.A_i(comb[9][9]), .B_i(comb[10][8]), .c_in(comb[11][7]), .S_o(S_s6_18_3), .c_out(C_s6_18_3));
logic S_s6_18_4, C_s6_18_4;
FA FA_s6_18_4(.A_i(comb[12][6]), .B_i(comb[13][5]), .c_in(comb[14][4]), .S_o(S_s6_18_4), .c_out(C_s6_18_4));
logic S_s6_18_5, C_s6_18_5;
HA HA_s6_185(.A_i(comb[15][3]), .B_i(comb[16][2]), .S_o(S_s6_18_5), .c_out(C_s6_18_5));
logic S_s6_19_0, C_s6_19_0;
FA FA_s6_19_0(.A_i(S_s7_19_0), .B_i(comb[2][17]), .c_in(comb[3][16]), .S_o(S_s6_19_0), .c_out(C_s6_19_0));
logic S_s6_19_1, C_s6_19_1;
FA FA_s6_19_1(.A_i(comb[4][15]), .B_i(comb[5][14]), .c_in(comb[6][13]), .S_o(S_s6_19_1), .c_out(C_s6_19_1));
logic S_s6_19_2, C_s6_19_2;
FA FA_s6_19_2(.A_i(comb[7][12]), .B_i(comb[8][11]), .c_in(comb[9][10]), .S_o(S_s6_19_2), .c_out(C_s6_19_2));
logic S_s6_19_3, C_s6_19_3;
FA FA_s6_19_3(.A_i(comb[10][9]), .B_i(comb[11][8]), .c_in(comb[12][7]), .S_o(S_s6_19_3), .c_out(C_s6_19_3));
logic S_s6_19_4, C_s6_19_4;
FA FA_s6_19_4(.A_i(comb[13][6]), .B_i(comb[14][5]), .c_in(comb[15][4]), .S_o(S_s6_19_4), .c_out(C_s6_19_4));
logic S_s6_19_5, C_s6_19_5;
FA FA_s6_19_5(.A_i(comb[16][3]), .B_i(comb[17][2]), .c_in(comb[18][1]), .S_o(S_s6_19_5), .c_out(C_s6_19_5));
logic S_s6_20_0, C_s6_20_0;
FA FA_s6_20_0(.A_i(S_s7_20_1), .B_i(S_s7_20_0), .c_in(C_s7_19_0), .S_o(S_s6_20_0), .c_out(C_s6_20_0));
logic S_s6_20_1, C_s6_20_1;
FA FA_s6_20_1(.A_i(comb[5][15]), .B_i(comb[6][14]), .c_in(comb[7][13]), .S_o(S_s6_20_1), .c_out(C_s6_20_1));
logic S_s6_20_2, C_s6_20_2;
FA FA_s6_20_2(.A_i(comb[8][12]), .B_i(comb[9][11]), .c_in(comb[10][10]), .S_o(S_s6_20_2), .c_out(C_s6_20_2));
logic S_s6_20_3, C_s6_20_3;
FA FA_s6_20_3(.A_i(comb[11][9]), .B_i(comb[12][8]), .c_in(comb[13][7]), .S_o(S_s6_20_3), .c_out(C_s6_20_3));
logic S_s6_20_4, C_s6_20_4;
FA FA_s6_20_4(.A_i(comb[14][6]), .B_i(comb[15][5]), .c_in(comb[16][4]), .S_o(S_s6_20_4), .c_out(C_s6_20_4));
logic S_s6_20_5, C_s6_20_5;
FA FA_s6_20_5(.A_i(comb[17][3]), .B_i(comb[18][2]), .c_in(comb[19][1]), .S_o(S_s6_20_5), .c_out(C_s6_20_5));
logic S_s6_21_0, C_s6_21_0;
FA FA_s6_21_0(.A_i(S_s7_21_2), .B_i(S_s7_21_1), .c_in(S_s7_21_0), .S_o(S_s6_21_0), .c_out(C_s6_21_0));
logic S_s6_21_1, C_s6_21_1;
FA FA_s6_21_1(.A_i(C_s7_20_1), .B_i(C_s7_20_0), .c_in(comb[8][13]), .S_o(S_s6_21_1), .c_out(C_s6_21_1));
logic S_s6_21_2, C_s6_21_2;
FA FA_s6_21_2(.A_i(comb[9][12]), .B_i(comb[10][11]), .c_in(comb[11][10]), .S_o(S_s6_21_2), .c_out(C_s6_21_2));
logic S_s6_21_3, C_s6_21_3;
FA FA_s6_21_3(.A_i(comb[12][9]), .B_i(comb[13][8]), .c_in(comb[14][7]), .S_o(S_s6_21_3), .c_out(C_s6_21_3));
logic S_s6_21_4, C_s6_21_4;
FA FA_s6_21_4(.A_i(comb[15][6]), .B_i(comb[16][5]), .c_in(comb[17][4]), .S_o(S_s6_21_4), .c_out(C_s6_21_4));
logic S_s6_21_5, C_s6_21_5;
FA FA_s6_21_5(.A_i(comb[18][3]), .B_i(comb[19][2]), .c_in(comb[20][1]), .S_o(S_s6_21_5), .c_out(C_s6_21_5));
logic S_s6_22_0, C_s6_22_0;
FA FA_s6_22_0(.A_i(S_s7_22_3), .B_i(S_s7_22_2), .c_in(S_s7_22_1), .S_o(S_s6_22_0), .c_out(C_s6_22_0));
logic S_s6_22_1, C_s6_22_1;
FA FA_s6_22_1(.A_i(S_s7_22_0), .B_i(C_s7_21_2), .c_in(C_s7_21_1), .S_o(S_s6_22_1), .c_out(C_s6_22_1));
logic S_s6_22_2, C_s6_22_2;
FA FA_s6_22_2(.A_i(C_s7_21_0), .B_i(comb[11][11]), .c_in(comb[12][10]), .S_o(S_s6_22_2), .c_out(C_s6_22_2));
logic S_s6_22_3, C_s6_22_3;
FA FA_s6_22_3(.A_i(comb[13][9]), .B_i(comb[14][8]), .c_in(comb[15][7]), .S_o(S_s6_22_3), .c_out(C_s6_22_3));
logic S_s6_22_4, C_s6_22_4;
FA FA_s6_22_4(.A_i(comb[16][6]), .B_i(comb[17][5]), .c_in(comb[18][4]), .S_o(S_s6_22_4), .c_out(C_s6_22_4));
logic S_s6_22_5, C_s6_22_5;
FA FA_s6_22_5(.A_i(comb[19][3]), .B_i(comb[20][2]), .c_in(comb[21][1]), .S_o(S_s6_22_5), .c_out(C_s6_22_5));
logic S_s6_23_0, C_s6_23_0;
FA FA_s6_23_0(.A_i(S_s7_23_4), .B_i(S_s7_23_3), .c_in(S_s7_23_2), .S_o(S_s6_23_0), .c_out(C_s6_23_0));
logic S_s6_23_1, C_s6_23_1;
FA FA_s6_23_1(.A_i(S_s7_23_1), .B_i(S_s7_23_0), .c_in(C_s7_22_3), .S_o(S_s6_23_1), .c_out(C_s6_23_1));
logic S_s6_23_2, C_s6_23_2;
FA FA_s6_23_2(.A_i(C_s7_22_2), .B_i(C_s7_22_1), .c_in(C_s7_22_0), .S_o(S_s6_23_2), .c_out(C_s6_23_2));
logic S_s6_23_3, C_s6_23_3;
FA FA_s6_23_3(.A_i(comb[14][9]), .B_i(comb[15][8]), .c_in(comb[16][7]), .S_o(S_s6_23_3), .c_out(C_s6_23_3));
logic S_s6_23_4, C_s6_23_4;
FA FA_s6_23_4(.A_i(comb[17][6]), .B_i(comb[18][5]), .c_in(comb[19][4]), .S_o(S_s6_23_4), .c_out(C_s6_23_4));
logic S_s6_23_5, C_s6_23_5;
FA FA_s6_23_5(.A_i(comb[20][3]), .B_i(comb[21][2]), .c_in(comb[22][1]), .S_o(S_s6_23_5), .c_out(C_s6_23_5));
logic S_s6_24_0, C_s6_24_0;
FA FA_s6_24_0(.A_i(S_s7_24_5), .B_i(S_s7_24_4), .c_in(S_s7_24_3), .S_o(S_s6_24_0), .c_out(C_s6_24_0));
logic S_s6_24_1, C_s6_24_1;
FA FA_s6_24_1(.A_i(S_s7_24_2), .B_i(S_s7_24_1), .c_in(S_s7_24_0), .S_o(S_s6_24_1), .c_out(C_s6_24_1));
logic S_s6_24_2, C_s6_24_2;
FA FA_s6_24_2(.A_i(C_s7_23_4), .B_i(C_s7_23_3), .c_in(C_s7_23_2), .S_o(S_s6_24_2), .c_out(C_s6_24_2));
logic S_s6_24_3, C_s6_24_3;
FA FA_s6_24_3(.A_i(C_s7_23_1), .B_i(C_s7_23_0), .c_in(comb[17][7]), .S_o(S_s6_24_3), .c_out(C_s6_24_3));
logic S_s6_24_4, C_s6_24_4;
FA FA_s6_24_4(.A_i(comb[18][6]), .B_i(comb[19][5]), .c_in(comb[20][4]), .S_o(S_s6_24_4), .c_out(C_s6_24_4));
logic S_s6_24_5, C_s6_24_5;
FA FA_s6_24_5(.A_i(comb[21][3]), .B_i(comb[22][2]), .c_in(comb[23][1]), .S_o(S_s6_24_5), .c_out(C_s6_24_5));
logic S_s6_25_0, C_s6_25_0;
FA FA_s6_25_0(.A_i(S_s7_25_6), .B_i(S_s7_25_5), .c_in(S_s7_25_4), .S_o(S_s6_25_0), .c_out(C_s6_25_0));
logic S_s6_25_1, C_s6_25_1;
FA FA_s6_25_1(.A_i(S_s7_25_3), .B_i(S_s7_25_2), .c_in(S_s7_25_1), .S_o(S_s6_25_1), .c_out(C_s6_25_1));
logic S_s6_25_2, C_s6_25_2;
FA FA_s6_25_2(.A_i(S_s7_25_0), .B_i(C_s7_24_5), .c_in(C_s7_24_4), .S_o(S_s6_25_2), .c_out(C_s6_25_2));
logic S_s6_25_3, C_s6_25_3;
FA FA_s6_25_3(.A_i(C_s7_24_3), .B_i(C_s7_24_2), .c_in(C_s7_24_1), .S_o(S_s6_25_3), .c_out(C_s6_25_3));
logic S_s6_25_4, C_s6_25_4;
FA FA_s6_25_4(.A_i(C_s7_24_0), .B_i(comb[20][5]), .c_in(comb[21][4]), .S_o(S_s6_25_4), .c_out(C_s6_25_4));
logic S_s6_25_5, C_s6_25_5;
FA FA_s6_25_5(.A_i(comb[22][3]), .B_i(comb[23][2]), .c_in(comb[24][1]), .S_o(S_s6_25_5), .c_out(C_s6_25_5));
logic S_s6_26_0, C_s6_26_0;
FA FA_s6_26_0(.A_i(S_s7_26_7), .B_i(S_s7_26_6), .c_in(S_s7_26_5), .S_o(S_s6_26_0), .c_out(C_s6_26_0));
logic S_s6_26_1, C_s6_26_1;
FA FA_s6_26_1(.A_i(S_s7_26_4), .B_i(S_s7_26_3), .c_in(S_s7_26_2), .S_o(S_s6_26_1), .c_out(C_s6_26_1));
logic S_s6_26_2, C_s6_26_2;
FA FA_s6_26_2(.A_i(S_s7_26_1), .B_i(S_s7_26_0), .c_in(C_s7_25_6), .S_o(S_s6_26_2), .c_out(C_s6_26_2));
logic S_s6_26_3, C_s6_26_3;
FA FA_s6_26_3(.A_i(C_s7_25_5), .B_i(C_s7_25_4), .c_in(C_s7_25_3), .S_o(S_s6_26_3), .c_out(C_s6_26_3));
logic S_s6_26_4, C_s6_26_4;
FA FA_s6_26_4(.A_i(C_s7_25_2), .B_i(C_s7_25_1), .c_in(C_s7_25_0), .S_o(S_s6_26_4), .c_out(C_s6_26_4));
logic S_s6_26_5, C_s6_26_5;
FA FA_s6_26_5(.A_i(comb[23][3]), .B_i(comb[24][2]), .c_in(comb[25][1]), .S_o(S_s6_26_5), .c_out(C_s6_26_5));
logic S_s6_27_0, C_s6_27_0;
FA FA_s6_27_0(.A_i(S_s7_27_8), .B_i(S_s7_27_7), .c_in(S_s7_27_6), .S_o(S_s6_27_0), .c_out(C_s6_27_0));
logic S_s6_27_1, C_s6_27_1;
FA FA_s6_27_1(.A_i(S_s7_27_5), .B_i(S_s7_27_4), .c_in(S_s7_27_3), .S_o(S_s6_27_1), .c_out(C_s6_27_1));
logic S_s6_27_2, C_s6_27_2;
FA FA_s6_27_2(.A_i(S_s7_27_2), .B_i(S_s7_27_1), .c_in(S_s7_27_0), .S_o(S_s6_27_2), .c_out(C_s6_27_2));
logic S_s6_27_3, C_s6_27_3;
FA FA_s6_27_3(.A_i(C_s7_26_7), .B_i(C_s7_26_6), .c_in(C_s7_26_5), .S_o(S_s6_27_3), .c_out(C_s6_27_3));
logic S_s6_27_4, C_s6_27_4;
FA FA_s6_27_4(.A_i(C_s7_26_4), .B_i(C_s7_26_3), .c_in(C_s7_26_2), .S_o(S_s6_27_4), .c_out(C_s6_27_4));
logic S_s6_27_5, C_s6_27_5;
FA FA_s6_27_5(.A_i(C_s7_26_1), .B_i(C_s7_26_0), .c_in(comb[26][1]), .S_o(S_s6_27_5), .c_out(C_s6_27_5));
logic S_s6_28_0, C_s6_28_0;
FA FA_s6_28_0(.A_i(S_s7_28_8), .B_i(S_s7_28_7), .c_in(S_s7_28_6), .S_o(S_s6_28_0), .c_out(C_s6_28_0));
logic S_s6_28_1, C_s6_28_1;
FA FA_s6_28_1(.A_i(S_s7_28_5), .B_i(S_s7_28_4), .c_in(S_s7_28_3), .S_o(S_s6_28_1), .c_out(C_s6_28_1));
logic S_s6_28_2, C_s6_28_2;
FA FA_s6_28_2(.A_i(S_s7_28_2), .B_i(S_s7_28_1), .c_in(S_s7_28_0), .S_o(S_s6_28_2), .c_out(C_s6_28_2));
logic S_s6_28_3, C_s6_28_3;
FA FA_s6_28_3(.A_i(C_s7_27_8), .B_i(C_s7_27_7), .c_in(C_s7_27_6), .S_o(S_s6_28_3), .c_out(C_s6_28_3));
logic S_s6_28_4, C_s6_28_4;
FA FA_s6_28_4(.A_i(C_s7_27_5), .B_i(C_s7_27_4), .c_in(C_s7_27_3), .S_o(S_s6_28_4), .c_out(C_s6_28_4));
logic S_s6_28_5, C_s6_28_5;
FA FA_s6_28_5(.A_i(C_s7_27_2), .B_i(C_s7_27_1), .c_in(C_s7_27_0), .S_o(S_s6_28_5), .c_out(C_s6_28_5));
logic S_s6_29_0, C_s6_29_0;
FA FA_s6_29_0(.A_i(S_s7_29_8), .B_i(S_s7_29_7), .c_in(S_s7_29_6), .S_o(S_s6_29_0), .c_out(C_s6_29_0));
logic S_s6_29_1, C_s6_29_1;
FA FA_s6_29_1(.A_i(S_s7_29_5), .B_i(S_s7_29_4), .c_in(S_s7_29_3), .S_o(S_s6_29_1), .c_out(C_s6_29_1));
logic S_s6_29_2, C_s6_29_2;
FA FA_s6_29_2(.A_i(S_s7_29_2), .B_i(S_s7_29_1), .c_in(S_s7_29_0), .S_o(S_s6_29_2), .c_out(C_s6_29_2));
logic S_s6_29_3, C_s6_29_3;
FA FA_s6_29_3(.A_i(C_s7_28_8), .B_i(C_s7_28_7), .c_in(C_s7_28_6), .S_o(S_s6_29_3), .c_out(C_s6_29_3));
logic S_s6_29_4, C_s6_29_4;
FA FA_s6_29_4(.A_i(C_s7_28_5), .B_i(C_s7_28_4), .c_in(C_s7_28_3), .S_o(S_s6_29_4), .c_out(C_s6_29_4));
logic S_s6_29_5, C_s6_29_5;
FA FA_s6_29_5(.A_i(C_s7_28_2), .B_i(C_s7_28_1), .c_in(C_s7_28_0), .S_o(S_s6_29_5), .c_out(C_s6_29_5));
logic S_s6_30_0, C_s6_30_0;
FA FA_s6_30_0(.A_i(S_s7_30_8), .B_i(S_s7_30_7), .c_in(S_s7_30_6), .S_o(S_s6_30_0), .c_out(C_s6_30_0));
logic S_s6_30_1, C_s6_30_1;
FA FA_s6_30_1(.A_i(S_s7_30_5), .B_i(S_s7_30_4), .c_in(S_s7_30_3), .S_o(S_s6_30_1), .c_out(C_s6_30_1));
logic S_s6_30_2, C_s6_30_2;
FA FA_s6_30_2(.A_i(S_s7_30_2), .B_i(S_s7_30_1), .c_in(S_s7_30_0), .S_o(S_s6_30_2), .c_out(C_s6_30_2));
logic S_s6_30_3, C_s6_30_3;
FA FA_s6_30_3(.A_i(C_s7_29_8), .B_i(C_s7_29_7), .c_in(C_s7_29_6), .S_o(S_s6_30_3), .c_out(C_s6_30_3));
logic S_s6_30_4, C_s6_30_4;
FA FA_s6_30_4(.A_i(C_s7_29_5), .B_i(C_s7_29_4), .c_in(C_s7_29_3), .S_o(S_s6_30_4), .c_out(C_s6_30_4));
logic S_s6_30_5, C_s6_30_5;
FA FA_s6_30_5(.A_i(C_s7_29_2), .B_i(C_s7_29_1), .c_in(C_s7_29_0), .S_o(S_s6_30_5), .c_out(C_s6_30_5));
logic S_s6_31_0, C_s6_31_0;
FA FA_s6_31_0(.A_i(S_s7_31_8), .B_i(S_s7_31_7), .c_in(S_s7_31_6), .S_o(S_s6_31_0), .c_out(C_s6_31_0));
logic S_s6_31_1, C_s6_31_1;
FA FA_s6_31_1(.A_i(S_s7_31_5), .B_i(S_s7_31_4), .c_in(S_s7_31_3), .S_o(S_s6_31_1), .c_out(C_s6_31_1));
logic S_s6_31_2, C_s6_31_2;
FA FA_s6_31_2(.A_i(S_s7_31_2), .B_i(S_s7_31_1), .c_in(S_s7_31_0), .S_o(S_s6_31_2), .c_out(C_s6_31_2));
logic S_s6_31_3, C_s6_31_3;
FA FA_s6_31_3(.A_i(C_s7_30_8), .B_i(C_s7_30_7), .c_in(C_s7_30_6), .S_o(S_s6_31_3), .c_out(C_s6_31_3));
logic S_s6_31_4, C_s6_31_4;
FA FA_s6_31_4(.A_i(C_s7_30_5), .B_i(C_s7_30_4), .c_in(C_s7_30_3), .S_o(S_s6_31_4), .c_out(C_s6_31_4));
logic S_s6_31_5, C_s6_31_5;
FA FA_s6_31_5(.A_i(C_s7_30_2), .B_i(C_s7_30_1), .c_in(C_s7_30_0), .S_o(S_s6_31_5), .c_out(C_s6_31_5));
logic S_s6_32_0, C_s6_32_0;
FA FA_s6_32_0(.A_i(S_s7_32_8), .B_i(S_s7_32_7), .c_in(S_s7_32_6), .S_o(S_s6_32_0), .c_out(C_s6_32_0));
logic S_s6_32_1, C_s6_32_1;
FA FA_s6_32_1(.A_i(S_s7_32_5), .B_i(S_s7_32_4), .c_in(S_s7_32_3), .S_o(S_s6_32_1), .c_out(C_s6_32_1));
logic S_s6_32_2, C_s6_32_2;
FA FA_s6_32_2(.A_i(S_s7_32_2), .B_i(S_s7_32_1), .c_in(S_s7_32_0), .S_o(S_s6_32_2), .c_out(C_s6_32_2));
logic S_s6_32_3, C_s6_32_3;
FA FA_s6_32_3(.A_i(C_s7_31_8), .B_i(C_s7_31_7), .c_in(C_s7_31_6), .S_o(S_s6_32_3), .c_out(C_s6_32_3));
logic S_s6_32_4, C_s6_32_4;
FA FA_s6_32_4(.A_i(C_s7_31_5), .B_i(C_s7_31_4), .c_in(C_s7_31_3), .S_o(S_s6_32_4), .c_out(C_s6_32_4));
logic S_s6_32_5, C_s6_32_5;
FA FA_s6_32_5(.A_i(C_s7_31_2), .B_i(C_s7_31_1), .c_in(C_s7_31_0), .S_o(S_s6_32_5), .c_out(C_s6_32_5));
logic S_s6_33_0, C_s6_33_0;
FA FA_s6_33_0(.A_i(S_s7_33_8), .B_i(S_s7_33_7), .c_in(S_s7_33_6), .S_o(S_s6_33_0), .c_out(C_s6_33_0));
logic S_s6_33_1, C_s6_33_1;
FA FA_s6_33_1(.A_i(S_s7_33_5), .B_i(S_s7_33_4), .c_in(S_s7_33_3), .S_o(S_s6_33_1), .c_out(C_s6_33_1));
logic S_s6_33_2, C_s6_33_2;
FA FA_s6_33_2(.A_i(S_s7_33_2), .B_i(S_s7_33_1), .c_in(S_s7_33_0), .S_o(S_s6_33_2), .c_out(C_s6_33_2));
logic S_s6_33_3, C_s6_33_3;
FA FA_s6_33_3(.A_i(C_s7_32_8), .B_i(C_s7_32_7), .c_in(C_s7_32_6), .S_o(S_s6_33_3), .c_out(C_s6_33_3));
logic S_s6_33_4, C_s6_33_4;
FA FA_s6_33_4(.A_i(C_s7_32_5), .B_i(C_s7_32_4), .c_in(C_s7_32_3), .S_o(S_s6_33_4), .c_out(C_s6_33_4));
logic S_s6_33_5, C_s6_33_5;
FA FA_s6_33_5(.A_i(C_s7_32_2), .B_i(C_s7_32_1), .c_in(C_s7_32_0), .S_o(S_s6_33_5), .c_out(C_s6_33_5));
logic S_s6_34_0, C_s6_34_0;
FA FA_s6_34_0(.A_i(S_s7_34_8), .B_i(S_s7_34_7), .c_in(S_s7_34_6), .S_o(S_s6_34_0), .c_out(C_s6_34_0));
logic S_s6_34_1, C_s6_34_1;
FA FA_s6_34_1(.A_i(S_s7_34_5), .B_i(S_s7_34_4), .c_in(S_s7_34_3), .S_o(S_s6_34_1), .c_out(C_s6_34_1));
logic S_s6_34_2, C_s6_34_2;
FA FA_s6_34_2(.A_i(S_s7_34_2), .B_i(S_s7_34_1), .c_in(S_s7_34_0), .S_o(S_s6_34_2), .c_out(C_s6_34_2));
logic S_s6_34_3, C_s6_34_3;
FA FA_s6_34_3(.A_i(C_s7_33_8), .B_i(C_s7_33_7), .c_in(C_s7_33_6), .S_o(S_s6_34_3), .c_out(C_s6_34_3));
logic S_s6_34_4, C_s6_34_4;
FA FA_s6_34_4(.A_i(C_s7_33_5), .B_i(C_s7_33_4), .c_in(C_s7_33_3), .S_o(S_s6_34_4), .c_out(C_s6_34_4));
logic S_s6_34_5, C_s6_34_5;
FA FA_s6_34_5(.A_i(C_s7_33_2), .B_i(C_s7_33_1), .c_in(C_s7_33_0), .S_o(S_s6_34_5), .c_out(C_s6_34_5));
logic S_s6_35_0, C_s6_35_0;
FA FA_s6_35_0(.A_i(S_s7_35_8), .B_i(S_s7_35_7), .c_in(S_s7_35_6), .S_o(S_s6_35_0), .c_out(C_s6_35_0));
logic S_s6_35_1, C_s6_35_1;
FA FA_s6_35_1(.A_i(S_s7_35_5), .B_i(S_s7_35_4), .c_in(S_s7_35_3), .S_o(S_s6_35_1), .c_out(C_s6_35_1));
logic S_s6_35_2, C_s6_35_2;
FA FA_s6_35_2(.A_i(S_s7_35_2), .B_i(S_s7_35_1), .c_in(S_s7_35_0), .S_o(S_s6_35_2), .c_out(C_s6_35_2));
logic S_s6_35_3, C_s6_35_3;
FA FA_s6_35_3(.A_i(C_s7_34_8), .B_i(C_s7_34_7), .c_in(C_s7_34_6), .S_o(S_s6_35_3), .c_out(C_s6_35_3));
logic S_s6_35_4, C_s6_35_4;
FA FA_s6_35_4(.A_i(C_s7_34_5), .B_i(C_s7_34_4), .c_in(C_s7_34_3), .S_o(S_s6_35_4), .c_out(C_s6_35_4));
logic S_s6_35_5, C_s6_35_5;
FA FA_s6_35_5(.A_i(C_s7_34_2), .B_i(C_s7_34_1), .c_in(C_s7_34_0), .S_o(S_s6_35_5), .c_out(C_s6_35_5));
logic S_s6_36_0, C_s6_36_0;
FA FA_s6_36_0(.A_i(S_s7_36_8), .B_i(S_s7_36_7), .c_in(S_s7_36_6), .S_o(S_s6_36_0), .c_out(C_s6_36_0));
logic S_s6_36_1, C_s6_36_1;
FA FA_s6_36_1(.A_i(S_s7_36_5), .B_i(S_s7_36_4), .c_in(S_s7_36_3), .S_o(S_s6_36_1), .c_out(C_s6_36_1));
logic S_s6_36_2, C_s6_36_2;
FA FA_s6_36_2(.A_i(S_s7_36_2), .B_i(S_s7_36_1), .c_in(S_s7_36_0), .S_o(S_s6_36_2), .c_out(C_s6_36_2));
logic S_s6_36_3, C_s6_36_3;
FA FA_s6_36_3(.A_i(C_s7_35_8), .B_i(C_s7_35_7), .c_in(C_s7_35_6), .S_o(S_s6_36_3), .c_out(C_s6_36_3));
logic S_s6_36_4, C_s6_36_4;
FA FA_s6_36_4(.A_i(C_s7_35_5), .B_i(C_s7_35_4), .c_in(C_s7_35_3), .S_o(S_s6_36_4), .c_out(C_s6_36_4));
logic S_s6_36_5, C_s6_36_5;
FA FA_s6_36_5(.A_i(C_s7_35_2), .B_i(C_s7_35_1), .c_in(C_s7_35_0), .S_o(S_s6_36_5), .c_out(C_s6_36_5));
logic S_s6_37_0, C_s6_37_0;
FA FA_s6_37_0(.A_i(S_s7_37_7), .B_i(S_s7_37_6), .c_in(S_s7_37_5), .S_o(S_s6_37_0), .c_out(C_s6_37_0));
logic S_s6_37_1, C_s6_37_1;
FA FA_s6_37_1(.A_i(S_s7_37_4), .B_i(S_s7_37_3), .c_in(S_s7_37_2), .S_o(S_s6_37_1), .c_out(C_s6_37_1));
logic S_s6_37_2, C_s6_37_2;
FA FA_s6_37_2(.A_i(S_s7_37_1), .B_i(S_s7_37_0), .c_in(C_s7_36_8), .S_o(S_s6_37_2), .c_out(C_s6_37_2));
logic S_s6_37_3, C_s6_37_3;
FA FA_s6_37_3(.A_i(C_s7_36_7), .B_i(C_s7_36_6), .c_in(C_s7_36_5), .S_o(S_s6_37_3), .c_out(C_s6_37_3));
logic S_s6_37_4, C_s6_37_4;
FA FA_s6_37_4(.A_i(C_s7_36_4), .B_i(C_s7_36_3), .c_in(C_s7_36_2), .S_o(S_s6_37_4), .c_out(C_s6_37_4));
logic S_s6_37_5, C_s6_37_5;
FA FA_s6_37_5(.A_i(C_s7_36_1), .B_i(C_s7_36_0), .c_in(comb[30][7]), .S_o(S_s6_37_5), .c_out(C_s6_37_5));
logic S_s6_38_0, C_s6_38_0;
FA FA_s6_38_0(.A_i(S_s7_38_6), .B_i(S_s7_38_5), .c_in(S_s7_38_4), .S_o(S_s6_38_0), .c_out(C_s6_38_0));
logic S_s6_38_1, C_s6_38_1;
FA FA_s6_38_1(.A_i(S_s7_38_3), .B_i(S_s7_38_2), .c_in(S_s7_38_1), .S_o(S_s6_38_1), .c_out(C_s6_38_1));
logic S_s6_38_2, C_s6_38_2;
FA FA_s6_38_2(.A_i(S_s7_38_0), .B_i(C_s7_37_7), .c_in(C_s7_37_6), .S_o(S_s6_38_2), .c_out(C_s6_38_2));
logic S_s6_38_3, C_s6_38_3;
FA FA_s6_38_3(.A_i(C_s7_37_5), .B_i(C_s7_37_4), .c_in(C_s7_37_3), .S_o(S_s6_38_3), .c_out(C_s6_38_3));
logic S_s6_38_4, C_s6_38_4;
FA FA_s6_38_4(.A_i(C_s7_37_2), .B_i(C_s7_37_1), .c_in(C_s7_37_0), .S_o(S_s6_38_4), .c_out(C_s6_38_4));
logic S_s6_38_5, C_s6_38_5;
FA FA_s6_38_5(.A_i(comb[28][10]), .B_i(comb[29][9]), .c_in(comb[30][8]), .S_o(S_s6_38_5), .c_out(C_s6_38_5));
logic S_s6_39_0, C_s6_39_0;
FA FA_s6_39_0(.A_i(S_s7_39_5), .B_i(S_s7_39_4), .c_in(S_s7_39_3), .S_o(S_s6_39_0), .c_out(C_s6_39_0));
logic S_s6_39_1, C_s6_39_1;
FA FA_s6_39_1(.A_i(S_s7_39_2), .B_i(S_s7_39_1), .c_in(S_s7_39_0), .S_o(S_s6_39_1), .c_out(C_s6_39_1));
logic S_s6_39_2, C_s6_39_2;
FA FA_s6_39_2(.A_i(C_s7_38_6), .B_i(C_s7_38_5), .c_in(C_s7_38_4), .S_o(S_s6_39_2), .c_out(C_s6_39_2));
logic S_s6_39_3, C_s6_39_3;
FA FA_s6_39_3(.A_i(C_s7_38_3), .B_i(C_s7_38_2), .c_in(C_s7_38_1), .S_o(S_s6_39_3), .c_out(C_s6_39_3));
logic S_s6_39_4, C_s6_39_4;
FA FA_s6_39_4(.A_i(C_s7_38_0), .B_i(comb[26][13]), .c_in(comb[27][12]), .S_o(S_s6_39_4), .c_out(C_s6_39_4));
logic S_s6_39_5, C_s6_39_5;
FA FA_s6_39_5(.A_i(comb[28][11]), .B_i(comb[29][10]), .c_in(comb[30][9]), .S_o(S_s6_39_5), .c_out(C_s6_39_5));
logic S_s6_40_0, C_s6_40_0;
FA FA_s6_40_0(.A_i(S_s7_40_4), .B_i(S_s7_40_3), .c_in(S_s7_40_2), .S_o(S_s6_40_0), .c_out(C_s6_40_0));
logic S_s6_40_1, C_s6_40_1;
FA FA_s6_40_1(.A_i(S_s7_40_1), .B_i(S_s7_40_0), .c_in(C_s7_39_5), .S_o(S_s6_40_1), .c_out(C_s6_40_1));
logic S_s6_40_2, C_s6_40_2;
FA FA_s6_40_2(.A_i(C_s7_39_4), .B_i(C_s7_39_3), .c_in(C_s7_39_2), .S_o(S_s6_40_2), .c_out(C_s6_40_2));
logic S_s6_40_3, C_s6_40_3;
FA FA_s6_40_3(.A_i(C_s7_39_1), .B_i(C_s7_39_0), .c_in(comb[24][16]), .S_o(S_s6_40_3), .c_out(C_s6_40_3));
logic S_s6_40_4, C_s6_40_4;
FA FA_s6_40_4(.A_i(comb[25][15]), .B_i(comb[26][14]), .c_in(comb[27][13]), .S_o(S_s6_40_4), .c_out(C_s6_40_4));
logic S_s6_40_5, C_s6_40_5;
FA FA_s6_40_5(.A_i(comb[28][12]), .B_i(comb[29][11]), .c_in(comb[30][10]), .S_o(S_s6_40_5), .c_out(C_s6_40_5));
logic S_s6_41_0, C_s6_41_0;
FA FA_s6_41_0(.A_i(S_s7_41_3), .B_i(S_s7_41_2), .c_in(S_s7_41_1), .S_o(S_s6_41_0), .c_out(C_s6_41_0));
logic S_s6_41_1, C_s6_41_1;
FA FA_s6_41_1(.A_i(S_s7_41_0), .B_i(C_s7_40_4), .c_in(C_s7_40_3), .S_o(S_s6_41_1), .c_out(C_s6_41_1));
logic S_s6_41_2, C_s6_41_2;
FA FA_s6_41_2(.A_i(C_s7_40_2), .B_i(C_s7_40_1), .c_in(C_s7_40_0), .S_o(S_s6_41_2), .c_out(C_s6_41_2));
logic S_s6_41_3, C_s6_41_3;
FA FA_s6_41_3(.A_i(comb[22][19]), .B_i(comb[23][18]), .c_in(comb[24][17]), .S_o(S_s6_41_3), .c_out(C_s6_41_3));
logic S_s6_41_4, C_s6_41_4;
FA FA_s6_41_4(.A_i(comb[25][16]), .B_i(comb[26][15]), .c_in(comb[27][14]), .S_o(S_s6_41_4), .c_out(C_s6_41_4));
logic S_s6_41_5, C_s6_41_5;
FA FA_s6_41_5(.A_i(comb[28][13]), .B_i(comb[29][12]), .c_in(comb[30][11]), .S_o(S_s6_41_5), .c_out(C_s6_41_5));
logic S_s6_42_0, C_s6_42_0;
FA FA_s6_42_0(.A_i(S_s7_42_2), .B_i(S_s7_42_1), .c_in(S_s7_42_0), .S_o(S_s6_42_0), .c_out(C_s6_42_0));
logic S_s6_42_1, C_s6_42_1;
FA FA_s6_42_1(.A_i(C_s7_41_3), .B_i(C_s7_41_2), .c_in(C_s7_41_1), .S_o(S_s6_42_1), .c_out(C_s6_42_1));
logic S_s6_42_2, C_s6_42_2;
FA FA_s6_42_2(.A_i(C_s7_41_0), .B_i(comb[20][22]), .c_in(comb[21][21]), .S_o(S_s6_42_2), .c_out(C_s6_42_2));
logic S_s6_42_3, C_s6_42_3;
FA FA_s6_42_3(.A_i(comb[22][20]), .B_i(comb[23][19]), .c_in(comb[24][18]), .S_o(S_s6_42_3), .c_out(C_s6_42_3));
logic S_s6_42_4, C_s6_42_4;
FA FA_s6_42_4(.A_i(comb[25][17]), .B_i(comb[26][16]), .c_in(comb[27][15]), .S_o(S_s6_42_4), .c_out(C_s6_42_4));
logic S_s6_42_5, C_s6_42_5;
FA FA_s6_42_5(.A_i(comb[28][14]), .B_i(comb[29][13]), .c_in(comb[30][12]), .S_o(S_s6_42_5), .c_out(C_s6_42_5));
logic S_s6_43_0, C_s6_43_0;
FA FA_s6_43_0(.A_i(S_s7_43_1), .B_i(S_s7_43_0), .c_in(C_s7_42_2), .S_o(S_s6_43_0), .c_out(C_s6_43_0));
logic S_s6_43_1, C_s6_43_1;
FA FA_s6_43_1(.A_i(C_s7_42_1), .B_i(C_s7_42_0), .c_in(comb[18][25]), .S_o(S_s6_43_1), .c_out(C_s6_43_1));
logic S_s6_43_2, C_s6_43_2;
FA FA_s6_43_2(.A_i(comb[19][24]), .B_i(comb[20][23]), .c_in(comb[21][22]), .S_o(S_s6_43_2), .c_out(C_s6_43_2));
logic S_s6_43_3, C_s6_43_3;
FA FA_s6_43_3(.A_i(comb[22][21]), .B_i(comb[23][20]), .c_in(comb[24][19]), .S_o(S_s6_43_3), .c_out(C_s6_43_3));
logic S_s6_43_4, C_s6_43_4;
FA FA_s6_43_4(.A_i(comb[25][18]), .B_i(comb[26][17]), .c_in(comb[27][16]), .S_o(S_s6_43_4), .c_out(C_s6_43_4));
logic S_s6_43_5, C_s6_43_5;
FA FA_s6_43_5(.A_i(comb[28][15]), .B_i(comb[29][14]), .c_in(comb[30][13]), .S_o(S_s6_43_5), .c_out(C_s6_43_5));
logic S_s6_44_0, C_s6_44_0;
FA FA_s6_44_0(.A_i(S_s7_44_0), .B_i(C_s7_43_1), .c_in(C_s7_43_0), .S_o(S_s6_44_0), .c_out(C_s6_44_0));
logic S_s6_44_1, C_s6_44_1;
FA FA_s6_44_1(.A_i(comb[16][28]), .B_i(comb[17][27]), .c_in(comb[18][26]), .S_o(S_s6_44_1), .c_out(C_s6_44_1));
logic S_s6_44_2, C_s6_44_2;
FA FA_s6_44_2(.A_i(comb[19][25]), .B_i(comb[20][24]), .c_in(comb[21][23]), .S_o(S_s6_44_2), .c_out(C_s6_44_2));
logic S_s6_44_3, C_s6_44_3;
FA FA_s6_44_3(.A_i(comb[22][22]), .B_i(comb[23][21]), .c_in(comb[24][20]), .S_o(S_s6_44_3), .c_out(C_s6_44_3));
logic S_s6_44_4, C_s6_44_4;
FA FA_s6_44_4(.A_i(comb[25][19]), .B_i(comb[26][18]), .c_in(comb[27][17]), .S_o(S_s6_44_4), .c_out(C_s6_44_4));
logic S_s6_44_5, C_s6_44_5;
FA FA_s6_44_5(.A_i(comb[28][16]), .B_i(comb[29][15]), .c_in(comb[30][14]), .S_o(S_s6_44_5), .c_out(C_s6_44_5));
logic S_s6_45_0, C_s6_45_0;
FA FA_s6_45_0(.A_i(C_s7_44_0), .B_i(comb[14][31]), .c_in(comb[15][30]), .S_o(S_s6_45_0), .c_out(C_s6_45_0));
logic S_s6_45_1, C_s6_45_1;
FA FA_s6_45_1(.A_i(comb[16][29]), .B_i(comb[17][28]), .c_in(comb[18][27]), .S_o(S_s6_45_1), .c_out(C_s6_45_1));
logic S_s6_45_2, C_s6_45_2;
FA FA_s6_45_2(.A_i(comb[19][26]), .B_i(comb[20][25]), .c_in(comb[21][24]), .S_o(S_s6_45_2), .c_out(C_s6_45_2));
logic S_s6_45_3, C_s6_45_3;
FA FA_s6_45_3(.A_i(comb[22][23]), .B_i(comb[23][22]), .c_in(comb[24][21]), .S_o(S_s6_45_3), .c_out(C_s6_45_3));
logic S_s6_45_4, C_s6_45_4;
FA FA_s6_45_4(.A_i(comb[25][20]), .B_i(comb[26][19]), .c_in(comb[27][18]), .S_o(S_s6_45_4), .c_out(C_s6_45_4));
logic S_s6_45_5, C_s6_45_5;
FA FA_s6_45_5(.A_i(comb[28][17]), .B_i(comb[29][16]), .c_in(comb[30][15]), .S_o(S_s6_45_5), .c_out(C_s6_45_5));
logic S_s6_46_0, C_s6_46_0;
FA FA_s6_46_0(.A_i(comb[15][31]), .B_i(comb[16][30]), .c_in(comb[17][29]), .S_o(S_s6_46_0), .c_out(C_s6_46_0));
logic S_s6_46_1, C_s6_46_1;
FA FA_s6_46_1(.A_i(comb[18][28]), .B_i(comb[19][27]), .c_in(comb[20][26]), .S_o(S_s6_46_1), .c_out(C_s6_46_1));
logic S_s6_46_2, C_s6_46_2;
FA FA_s6_46_2(.A_i(comb[21][25]), .B_i(comb[22][24]), .c_in(comb[23][23]), .S_o(S_s6_46_2), .c_out(C_s6_46_2));
logic S_s6_46_3, C_s6_46_3;
FA FA_s6_46_3(.A_i(comb[24][22]), .B_i(comb[25][21]), .c_in(comb[26][20]), .S_o(S_s6_46_3), .c_out(C_s6_46_3));
logic S_s6_46_4, C_s6_46_4;
FA FA_s6_46_4(.A_i(comb[27][19]), .B_i(comb[28][18]), .c_in(comb[29][17]), .S_o(S_s6_46_4), .c_out(C_s6_46_4));
logic S_s6_47_0, C_s6_47_0;
FA FA_s6_47_0(.A_i(comb[16][31]), .B_i(comb[17][30]), .c_in(comb[18][29]), .S_o(S_s6_47_0), .c_out(C_s6_47_0));
logic S_s6_47_1, C_s6_47_1;
FA FA_s6_47_1(.A_i(comb[19][28]), .B_i(comb[20][27]), .c_in(comb[21][26]), .S_o(S_s6_47_1), .c_out(C_s6_47_1));
logic S_s6_47_2, C_s6_47_2;
FA FA_s6_47_2(.A_i(comb[22][25]), .B_i(comb[23][24]), .c_in(comb[24][23]), .S_o(S_s6_47_2), .c_out(C_s6_47_2));
logic S_s6_47_3, C_s6_47_3;
FA FA_s6_47_3(.A_i(comb[25][22]), .B_i(comb[26][21]), .c_in(comb[27][20]), .S_o(S_s6_47_3), .c_out(C_s6_47_3));
logic S_s6_48_0, C_s6_48_0;
FA FA_s6_48_0(.A_i(comb[17][31]), .B_i(comb[18][30]), .c_in(comb[19][29]), .S_o(S_s6_48_0), .c_out(C_s6_48_0));
logic S_s6_48_1, C_s6_48_1;
FA FA_s6_48_1(.A_i(comb[20][28]), .B_i(comb[21][27]), .c_in(comb[22][26]), .S_o(S_s6_48_1), .c_out(C_s6_48_1));
logic S_s6_48_2, C_s6_48_2;
FA FA_s6_48_2(.A_i(comb[23][25]), .B_i(comb[24][24]), .c_in(comb[25][23]), .S_o(S_s6_48_2), .c_out(C_s6_48_2));
logic S_s6_49_0, C_s6_49_0;
FA FA_s6_49_0(.A_i(comb[18][31]), .B_i(comb[19][30]), .c_in(comb[20][29]), .S_o(S_s6_49_0), .c_out(C_s6_49_0));
logic S_s6_49_1, C_s6_49_1;
FA FA_s6_49_1(.A_i(comb[21][28]), .B_i(comb[22][27]), .c_in(comb[23][26]), .S_o(S_s6_49_1), .c_out(C_s6_49_1));
logic S_s6_50_0, C_s6_50_0;
FA FA_s6_50_0(.A_i(comb[19][31]), .B_i(comb[20][30]), .c_in(comb[21][29]), .S_o(S_s6_50_0), .c_out(C_s6_50_0));
// stage 6 end ======================================================================================================= 

// stage 5 begin ======================================================================================================= 
logic S_s5_9_0, C_s5_9_0;
HA HA_s5_90(.A_i(comb[0][9]), .B_i(comb[1][8]), .S_o(S_s5_9_0), .c_out(C_s5_9_0));
logic S_s5_10_0, C_s5_10_0;
FA FA_s5_10_0(.A_i(comb[0][10]), .B_i(comb[1][9]), .c_in(comb[2][8]), .S_o(S_s5_10_0), .c_out(C_s5_10_0));
logic S_s5_10_1, C_s5_10_1;
HA HA_s5_101(.A_i(comb[3][7]), .B_i(comb[4][6]), .S_o(S_s5_10_1), .c_out(C_s5_10_1));
logic S_s5_11_0, C_s5_11_0;
FA FA_s5_11_0(.A_i(comb[0][11]), .B_i(comb[1][10]), .c_in(comb[2][9]), .S_o(S_s5_11_0), .c_out(C_s5_11_0));
logic S_s5_11_1, C_s5_11_1;
FA FA_s5_11_1(.A_i(comb[3][8]), .B_i(comb[4][7]), .c_in(comb[5][6]), .S_o(S_s5_11_1), .c_out(C_s5_11_1));
logic S_s5_11_2, C_s5_11_2;
HA HA_s5_112(.A_i(comb[6][5]), .B_i(comb[7][4]), .S_o(S_s5_11_2), .c_out(C_s5_11_2));
logic S_s5_12_0, C_s5_12_0;
FA FA_s5_12_0(.A_i(comb[0][12]), .B_i(comb[1][11]), .c_in(comb[2][10]), .S_o(S_s5_12_0), .c_out(C_s5_12_0));
logic S_s5_12_1, C_s5_12_1;
FA FA_s5_12_1(.A_i(comb[3][9]), .B_i(comb[4][8]), .c_in(comb[5][7]), .S_o(S_s5_12_1), .c_out(C_s5_12_1));
logic S_s5_12_2, C_s5_12_2;
FA FA_s5_12_2(.A_i(comb[6][6]), .B_i(comb[7][5]), .c_in(comb[8][4]), .S_o(S_s5_12_2), .c_out(C_s5_12_2));
logic S_s5_12_3, C_s5_12_3;
HA HA_s5_123(.A_i(comb[9][3]), .B_i(comb[10][2]), .S_o(S_s5_12_3), .c_out(C_s5_12_3));
logic S_s5_13_0, C_s5_13_0;
FA FA_s5_13_0(.A_i(S_s6_13_0), .B_i(comb[2][11]), .c_in(comb[3][10]), .S_o(S_s5_13_0), .c_out(C_s5_13_0));
logic S_s5_13_1, C_s5_13_1;
FA FA_s5_13_1(.A_i(comb[4][9]), .B_i(comb[5][8]), .c_in(comb[6][7]), .S_o(S_s5_13_1), .c_out(C_s5_13_1));
logic S_s5_13_2, C_s5_13_2;
FA FA_s5_13_2(.A_i(comb[7][6]), .B_i(comb[8][5]), .c_in(comb[9][4]), .S_o(S_s5_13_2), .c_out(C_s5_13_2));
logic S_s5_13_3, C_s5_13_3;
FA FA_s5_13_3(.A_i(comb[10][3]), .B_i(comb[11][2]), .c_in(comb[12][1]), .S_o(S_s5_13_3), .c_out(C_s5_13_3));
logic S_s5_14_0, C_s5_14_0;
FA FA_s5_14_0(.A_i(S_s6_14_1), .B_i(S_s6_14_0), .c_in(C_s6_13_0), .S_o(S_s5_14_0), .c_out(C_s5_14_0));
logic S_s5_14_1, C_s5_14_1;
FA FA_s5_14_1(.A_i(comb[5][9]), .B_i(comb[6][8]), .c_in(comb[7][7]), .S_o(S_s5_14_1), .c_out(C_s5_14_1));
logic S_s5_14_2, C_s5_14_2;
FA FA_s5_14_2(.A_i(comb[8][6]), .B_i(comb[9][5]), .c_in(comb[10][4]), .S_o(S_s5_14_2), .c_out(C_s5_14_2));
logic S_s5_14_3, C_s5_14_3;
FA FA_s5_14_3(.A_i(comb[11][3]), .B_i(comb[12][2]), .c_in(comb[13][1]), .S_o(S_s5_14_3), .c_out(C_s5_14_3));
logic S_s5_15_0, C_s5_15_0;
FA FA_s5_15_0(.A_i(S_s6_15_2), .B_i(S_s6_15_1), .c_in(S_s6_15_0), .S_o(S_s5_15_0), .c_out(C_s5_15_0));
logic S_s5_15_1, C_s5_15_1;
FA FA_s5_15_1(.A_i(C_s6_14_1), .B_i(C_s6_14_0), .c_in(comb[8][7]), .S_o(S_s5_15_1), .c_out(C_s5_15_1));
logic S_s5_15_2, C_s5_15_2;
FA FA_s5_15_2(.A_i(comb[9][6]), .B_i(comb[10][5]), .c_in(comb[11][4]), .S_o(S_s5_15_2), .c_out(C_s5_15_2));
logic S_s5_15_3, C_s5_15_3;
FA FA_s5_15_3(.A_i(comb[12][3]), .B_i(comb[13][2]), .c_in(comb[14][1]), .S_o(S_s5_15_3), .c_out(C_s5_15_3));
logic S_s5_16_0, C_s5_16_0;
FA FA_s5_16_0(.A_i(S_s6_16_3), .B_i(S_s6_16_2), .c_in(S_s6_16_1), .S_o(S_s5_16_0), .c_out(C_s5_16_0));
logic S_s5_16_1, C_s5_16_1;
FA FA_s5_16_1(.A_i(S_s6_16_0), .B_i(C_s6_15_2), .c_in(C_s6_15_1), .S_o(S_s5_16_1), .c_out(C_s5_16_1));
logic S_s5_16_2, C_s5_16_2;
FA FA_s5_16_2(.A_i(C_s6_15_0), .B_i(comb[11][5]), .c_in(comb[12][4]), .S_o(S_s5_16_2), .c_out(C_s5_16_2));
logic S_s5_16_3, C_s5_16_3;
FA FA_s5_16_3(.A_i(comb[13][3]), .B_i(comb[14][2]), .c_in(comb[15][1]), .S_o(S_s5_16_3), .c_out(C_s5_16_3));
logic S_s5_17_0, C_s5_17_0;
FA FA_s5_17_0(.A_i(S_s6_17_4), .B_i(S_s6_17_3), .c_in(S_s6_17_2), .S_o(S_s5_17_0), .c_out(C_s5_17_0));
logic S_s5_17_1, C_s5_17_1;
FA FA_s5_17_1(.A_i(S_s6_17_1), .B_i(S_s6_17_0), .c_in(C_s6_16_3), .S_o(S_s5_17_1), .c_out(C_s5_17_1));
logic S_s5_17_2, C_s5_17_2;
FA FA_s5_17_2(.A_i(C_s6_16_2), .B_i(C_s6_16_1), .c_in(C_s6_16_0), .S_o(S_s5_17_2), .c_out(C_s5_17_2));
logic S_s5_17_3, C_s5_17_3;
FA FA_s5_17_3(.A_i(comb[14][3]), .B_i(comb[15][2]), .c_in(comb[16][1]), .S_o(S_s5_17_3), .c_out(C_s5_17_3));
logic S_s5_18_0, C_s5_18_0;
FA FA_s5_18_0(.A_i(S_s6_18_5), .B_i(S_s6_18_4), .c_in(S_s6_18_3), .S_o(S_s5_18_0), .c_out(C_s5_18_0));
logic S_s5_18_1, C_s5_18_1;
FA FA_s5_18_1(.A_i(S_s6_18_2), .B_i(S_s6_18_1), .c_in(S_s6_18_0), .S_o(S_s5_18_1), .c_out(C_s5_18_1));
logic S_s5_18_2, C_s5_18_2;
FA FA_s5_18_2(.A_i(C_s6_17_4), .B_i(C_s6_17_3), .c_in(C_s6_17_2), .S_o(S_s5_18_2), .c_out(C_s5_18_2));
logic S_s5_18_3, C_s5_18_3;
FA FA_s5_18_3(.A_i(C_s6_17_1), .B_i(C_s6_17_0), .c_in(comb[17][1]), .S_o(S_s5_18_3), .c_out(C_s5_18_3));
logic S_s5_19_0, C_s5_19_0;
FA FA_s5_19_0(.A_i(S_s6_19_5), .B_i(S_s6_19_4), .c_in(S_s6_19_3), .S_o(S_s5_19_0), .c_out(C_s5_19_0));
logic S_s5_19_1, C_s5_19_1;
FA FA_s5_19_1(.A_i(S_s6_19_2), .B_i(S_s6_19_1), .c_in(S_s6_19_0), .S_o(S_s5_19_1), .c_out(C_s5_19_1));
logic S_s5_19_2, C_s5_19_2;
FA FA_s5_19_2(.A_i(C_s6_18_5), .B_i(C_s6_18_4), .c_in(C_s6_18_3), .S_o(S_s5_19_2), .c_out(C_s5_19_2));
logic S_s5_19_3, C_s5_19_3;
FA FA_s5_19_3(.A_i(C_s6_18_2), .B_i(C_s6_18_1), .c_in(C_s6_18_0), .S_o(S_s5_19_3), .c_out(C_s5_19_3));
logic S_s5_20_0, C_s5_20_0;
FA FA_s5_20_0(.A_i(S_s6_20_5), .B_i(S_s6_20_4), .c_in(S_s6_20_3), .S_o(S_s5_20_0), .c_out(C_s5_20_0));
logic S_s5_20_1, C_s5_20_1;
FA FA_s5_20_1(.A_i(S_s6_20_2), .B_i(S_s6_20_1), .c_in(S_s6_20_0), .S_o(S_s5_20_1), .c_out(C_s5_20_1));
logic S_s5_20_2, C_s5_20_2;
FA FA_s5_20_2(.A_i(C_s6_19_5), .B_i(C_s6_19_4), .c_in(C_s6_19_3), .S_o(S_s5_20_2), .c_out(C_s5_20_2));
logic S_s5_20_3, C_s5_20_3;
FA FA_s5_20_3(.A_i(C_s6_19_2), .B_i(C_s6_19_1), .c_in(C_s6_19_0), .S_o(S_s5_20_3), .c_out(C_s5_20_3));
logic S_s5_21_0, C_s5_21_0;
FA FA_s5_21_0(.A_i(S_s6_21_5), .B_i(S_s6_21_4), .c_in(S_s6_21_3), .S_o(S_s5_21_0), .c_out(C_s5_21_0));
logic S_s5_21_1, C_s5_21_1;
FA FA_s5_21_1(.A_i(S_s6_21_2), .B_i(S_s6_21_1), .c_in(S_s6_21_0), .S_o(S_s5_21_1), .c_out(C_s5_21_1));
logic S_s5_21_2, C_s5_21_2;
FA FA_s5_21_2(.A_i(C_s6_20_5), .B_i(C_s6_20_4), .c_in(C_s6_20_3), .S_o(S_s5_21_2), .c_out(C_s5_21_2));
logic S_s5_21_3, C_s5_21_3;
FA FA_s5_21_3(.A_i(C_s6_20_2), .B_i(C_s6_20_1), .c_in(C_s6_20_0), .S_o(S_s5_21_3), .c_out(C_s5_21_3));
logic S_s5_22_0, C_s5_22_0;
FA FA_s5_22_0(.A_i(S_s6_22_5), .B_i(S_s6_22_4), .c_in(S_s6_22_3), .S_o(S_s5_22_0), .c_out(C_s5_22_0));
logic S_s5_22_1, C_s5_22_1;
FA FA_s5_22_1(.A_i(S_s6_22_2), .B_i(S_s6_22_1), .c_in(S_s6_22_0), .S_o(S_s5_22_1), .c_out(C_s5_22_1));
logic S_s5_22_2, C_s5_22_2;
FA FA_s5_22_2(.A_i(C_s6_21_5), .B_i(C_s6_21_4), .c_in(C_s6_21_3), .S_o(S_s5_22_2), .c_out(C_s5_22_2));
logic S_s5_22_3, C_s5_22_3;
FA FA_s5_22_3(.A_i(C_s6_21_2), .B_i(C_s6_21_1), .c_in(C_s6_21_0), .S_o(S_s5_22_3), .c_out(C_s5_22_3));
logic S_s5_23_0, C_s5_23_0;
FA FA_s5_23_0(.A_i(S_s6_23_5), .B_i(S_s6_23_4), .c_in(S_s6_23_3), .S_o(S_s5_23_0), .c_out(C_s5_23_0));
logic S_s5_23_1, C_s5_23_1;
FA FA_s5_23_1(.A_i(S_s6_23_2), .B_i(S_s6_23_1), .c_in(S_s6_23_0), .S_o(S_s5_23_1), .c_out(C_s5_23_1));
logic S_s5_23_2, C_s5_23_2;
FA FA_s5_23_2(.A_i(C_s6_22_5), .B_i(C_s6_22_4), .c_in(C_s6_22_3), .S_o(S_s5_23_2), .c_out(C_s5_23_2));
logic S_s5_23_3, C_s5_23_3;
FA FA_s5_23_3(.A_i(C_s6_22_2), .B_i(C_s6_22_1), .c_in(C_s6_22_0), .S_o(S_s5_23_3), .c_out(C_s5_23_3));
logic S_s5_24_0, C_s5_24_0;
FA FA_s5_24_0(.A_i(S_s6_24_5), .B_i(S_s6_24_4), .c_in(S_s6_24_3), .S_o(S_s5_24_0), .c_out(C_s5_24_0));
logic S_s5_24_1, C_s5_24_1;
FA FA_s5_24_1(.A_i(S_s6_24_2), .B_i(S_s6_24_1), .c_in(S_s6_24_0), .S_o(S_s5_24_1), .c_out(C_s5_24_1));
logic S_s5_24_2, C_s5_24_2;
FA FA_s5_24_2(.A_i(C_s6_23_5), .B_i(C_s6_23_4), .c_in(C_s6_23_3), .S_o(S_s5_24_2), .c_out(C_s5_24_2));
logic S_s5_24_3, C_s5_24_3;
FA FA_s5_24_3(.A_i(C_s6_23_2), .B_i(C_s6_23_1), .c_in(C_s6_23_0), .S_o(S_s5_24_3), .c_out(C_s5_24_3));
logic S_s5_25_0, C_s5_25_0;
FA FA_s5_25_0(.A_i(S_s6_25_5), .B_i(S_s6_25_4), .c_in(S_s6_25_3), .S_o(S_s5_25_0), .c_out(C_s5_25_0));
logic S_s5_25_1, C_s5_25_1;
FA FA_s5_25_1(.A_i(S_s6_25_2), .B_i(S_s6_25_1), .c_in(S_s6_25_0), .S_o(S_s5_25_1), .c_out(C_s5_25_1));
logic S_s5_25_2, C_s5_25_2;
FA FA_s5_25_2(.A_i(C_s6_24_5), .B_i(C_s6_24_4), .c_in(C_s6_24_3), .S_o(S_s5_25_2), .c_out(C_s5_25_2));
logic S_s5_25_3, C_s5_25_3;
FA FA_s5_25_3(.A_i(C_s6_24_2), .B_i(C_s6_24_1), .c_in(C_s6_24_0), .S_o(S_s5_25_3), .c_out(C_s5_25_3));
logic S_s5_26_0, C_s5_26_0;
FA FA_s5_26_0(.A_i(S_s6_26_5), .B_i(S_s6_26_4), .c_in(S_s6_26_3), .S_o(S_s5_26_0), .c_out(C_s5_26_0));
logic S_s5_26_1, C_s5_26_1;
FA FA_s5_26_1(.A_i(S_s6_26_2), .B_i(S_s6_26_1), .c_in(S_s6_26_0), .S_o(S_s5_26_1), .c_out(C_s5_26_1));
logic S_s5_26_2, C_s5_26_2;
FA FA_s5_26_2(.A_i(C_s6_25_5), .B_i(C_s6_25_4), .c_in(C_s6_25_3), .S_o(S_s5_26_2), .c_out(C_s5_26_2));
logic S_s5_26_3, C_s5_26_3;
FA FA_s5_26_3(.A_i(C_s6_25_2), .B_i(C_s6_25_1), .c_in(C_s6_25_0), .S_o(S_s5_26_3), .c_out(C_s5_26_3));
logic S_s5_27_0, C_s5_27_0;
FA FA_s5_27_0(.A_i(S_s6_27_5), .B_i(S_s6_27_4), .c_in(S_s6_27_3), .S_o(S_s5_27_0), .c_out(C_s5_27_0));
logic S_s5_27_1, C_s5_27_1;
FA FA_s5_27_1(.A_i(S_s6_27_2), .B_i(S_s6_27_1), .c_in(S_s6_27_0), .S_o(S_s5_27_1), .c_out(C_s5_27_1));
logic S_s5_27_2, C_s5_27_2;
FA FA_s5_27_2(.A_i(C_s6_26_5), .B_i(C_s6_26_4), .c_in(C_s6_26_3), .S_o(S_s5_27_2), .c_out(C_s5_27_2));
logic S_s5_27_3, C_s5_27_3;
FA FA_s5_27_3(.A_i(C_s6_26_2), .B_i(C_s6_26_1), .c_in(C_s6_26_0), .S_o(S_s5_27_3), .c_out(C_s5_27_3));
logic S_s5_28_0, C_s5_28_0;
FA FA_s5_28_0(.A_i(S_s6_28_5), .B_i(S_s6_28_4), .c_in(S_s6_28_3), .S_o(S_s5_28_0), .c_out(C_s5_28_0));
logic S_s5_28_1, C_s5_28_1;
FA FA_s5_28_1(.A_i(S_s6_28_2), .B_i(S_s6_28_1), .c_in(S_s6_28_0), .S_o(S_s5_28_1), .c_out(C_s5_28_1));
logic S_s5_28_2, C_s5_28_2;
FA FA_s5_28_2(.A_i(C_s6_27_5), .B_i(C_s6_27_4), .c_in(C_s6_27_3), .S_o(S_s5_28_2), .c_out(C_s5_28_2));
logic S_s5_28_3, C_s5_28_3;
FA FA_s5_28_3(.A_i(C_s6_27_2), .B_i(C_s6_27_1), .c_in(C_s6_27_0), .S_o(S_s5_28_3), .c_out(C_s5_28_3));
logic S_s5_29_0, C_s5_29_0;
FA FA_s5_29_0(.A_i(S_s6_29_5), .B_i(S_s6_29_4), .c_in(S_s6_29_3), .S_o(S_s5_29_0), .c_out(C_s5_29_0));
logic S_s5_29_1, C_s5_29_1;
FA FA_s5_29_1(.A_i(S_s6_29_2), .B_i(S_s6_29_1), .c_in(S_s6_29_0), .S_o(S_s5_29_1), .c_out(C_s5_29_1));
logic S_s5_29_2, C_s5_29_2;
FA FA_s5_29_2(.A_i(C_s6_28_5), .B_i(C_s6_28_4), .c_in(C_s6_28_3), .S_o(S_s5_29_2), .c_out(C_s5_29_2));
logic S_s5_29_3, C_s5_29_3;
FA FA_s5_29_3(.A_i(C_s6_28_2), .B_i(C_s6_28_1), .c_in(C_s6_28_0), .S_o(S_s5_29_3), .c_out(C_s5_29_3));
logic S_s5_30_0, C_s5_30_0;
FA FA_s5_30_0(.A_i(S_s6_30_5), .B_i(S_s6_30_4), .c_in(S_s6_30_3), .S_o(S_s5_30_0), .c_out(C_s5_30_0));
logic S_s5_30_1, C_s5_30_1;
FA FA_s5_30_1(.A_i(S_s6_30_2), .B_i(S_s6_30_1), .c_in(S_s6_30_0), .S_o(S_s5_30_1), .c_out(C_s5_30_1));
logic S_s5_30_2, C_s5_30_2;
FA FA_s5_30_2(.A_i(C_s6_29_5), .B_i(C_s6_29_4), .c_in(C_s6_29_3), .S_o(S_s5_30_2), .c_out(C_s5_30_2));
logic S_s5_30_3, C_s5_30_3;
FA FA_s5_30_3(.A_i(C_s6_29_2), .B_i(C_s6_29_1), .c_in(C_s6_29_0), .S_o(S_s5_30_3), .c_out(C_s5_30_3));
logic S_s5_31_0, C_s5_31_0;
FA FA_s5_31_0(.A_i(S_s6_31_5), .B_i(S_s6_31_4), .c_in(S_s6_31_3), .S_o(S_s5_31_0), .c_out(C_s5_31_0));
logic S_s5_31_1, C_s5_31_1;
FA FA_s5_31_1(.A_i(S_s6_31_2), .B_i(S_s6_31_1), .c_in(S_s6_31_0), .S_o(S_s5_31_1), .c_out(C_s5_31_1));
logic S_s5_31_2, C_s5_31_2;
FA FA_s5_31_2(.A_i(C_s6_30_5), .B_i(C_s6_30_4), .c_in(C_s6_30_3), .S_o(S_s5_31_2), .c_out(C_s5_31_2));
logic S_s5_31_3, C_s5_31_3;
FA FA_s5_31_3(.A_i(C_s6_30_2), .B_i(C_s6_30_1), .c_in(C_s6_30_0), .S_o(S_s5_31_3), .c_out(C_s5_31_3));
logic S_s5_32_0, C_s5_32_0;
FA FA_s5_32_0(.A_i(S_s6_32_5), .B_i(S_s6_32_4), .c_in(S_s6_32_3), .S_o(S_s5_32_0), .c_out(C_s5_32_0));
logic S_s5_32_1, C_s5_32_1;
FA FA_s5_32_1(.A_i(S_s6_32_2), .B_i(S_s6_32_1), .c_in(S_s6_32_0), .S_o(S_s5_32_1), .c_out(C_s5_32_1));
logic S_s5_32_2, C_s5_32_2;
FA FA_s5_32_2(.A_i(C_s6_31_5), .B_i(C_s6_31_4), .c_in(C_s6_31_3), .S_o(S_s5_32_2), .c_out(C_s5_32_2));
logic S_s5_32_3, C_s5_32_3;
FA FA_s5_32_3(.A_i(C_s6_31_2), .B_i(C_s6_31_1), .c_in(C_s6_31_0), .S_o(S_s5_32_3), .c_out(C_s5_32_3));
logic S_s5_33_0, C_s5_33_0;
FA FA_s5_33_0(.A_i(S_s6_33_5), .B_i(S_s6_33_4), .c_in(S_s6_33_3), .S_o(S_s5_33_0), .c_out(C_s5_33_0));
logic S_s5_33_1, C_s5_33_1;
FA FA_s5_33_1(.A_i(S_s6_33_2), .B_i(S_s6_33_1), .c_in(S_s6_33_0), .S_o(S_s5_33_1), .c_out(C_s5_33_1));
logic S_s5_33_2, C_s5_33_2;
FA FA_s5_33_2(.A_i(C_s6_32_5), .B_i(C_s6_32_4), .c_in(C_s6_32_3), .S_o(S_s5_33_2), .c_out(C_s5_33_2));
logic S_s5_33_3, C_s5_33_3;
FA FA_s5_33_3(.A_i(C_s6_32_2), .B_i(C_s6_32_1), .c_in(C_s6_32_0), .S_o(S_s5_33_3), .c_out(C_s5_33_3));
logic S_s5_34_0, C_s5_34_0;
FA FA_s5_34_0(.A_i(S_s6_34_5), .B_i(S_s6_34_4), .c_in(S_s6_34_3), .S_o(S_s5_34_0), .c_out(C_s5_34_0));
logic S_s5_34_1, C_s5_34_1;
FA FA_s5_34_1(.A_i(S_s6_34_2), .B_i(S_s6_34_1), .c_in(S_s6_34_0), .S_o(S_s5_34_1), .c_out(C_s5_34_1));
logic S_s5_34_2, C_s5_34_2;
FA FA_s5_34_2(.A_i(C_s6_33_5), .B_i(C_s6_33_4), .c_in(C_s6_33_3), .S_o(S_s5_34_2), .c_out(C_s5_34_2));
logic S_s5_34_3, C_s5_34_3;
FA FA_s5_34_3(.A_i(C_s6_33_2), .B_i(C_s6_33_1), .c_in(C_s6_33_0), .S_o(S_s5_34_3), .c_out(C_s5_34_3));
logic S_s5_35_0, C_s5_35_0;
FA FA_s5_35_0(.A_i(S_s6_35_5), .B_i(S_s6_35_4), .c_in(S_s6_35_3), .S_o(S_s5_35_0), .c_out(C_s5_35_0));
logic S_s5_35_1, C_s5_35_1;
FA FA_s5_35_1(.A_i(S_s6_35_2), .B_i(S_s6_35_1), .c_in(S_s6_35_0), .S_o(S_s5_35_1), .c_out(C_s5_35_1));
logic S_s5_35_2, C_s5_35_2;
FA FA_s5_35_2(.A_i(C_s6_34_5), .B_i(C_s6_34_4), .c_in(C_s6_34_3), .S_o(S_s5_35_2), .c_out(C_s5_35_2));
logic S_s5_35_3, C_s5_35_3;
FA FA_s5_35_3(.A_i(C_s6_34_2), .B_i(C_s6_34_1), .c_in(C_s6_34_0), .S_o(S_s5_35_3), .c_out(C_s5_35_3));
logic S_s5_36_0, C_s5_36_0;
FA FA_s5_36_0(.A_i(S_s6_36_5), .B_i(S_s6_36_4), .c_in(S_s6_36_3), .S_o(S_s5_36_0), .c_out(C_s5_36_0));
logic S_s5_36_1, C_s5_36_1;
FA FA_s5_36_1(.A_i(S_s6_36_2), .B_i(S_s6_36_1), .c_in(S_s6_36_0), .S_o(S_s5_36_1), .c_out(C_s5_36_1));
logic S_s5_36_2, C_s5_36_2;
FA FA_s5_36_2(.A_i(C_s6_35_5), .B_i(C_s6_35_4), .c_in(C_s6_35_3), .S_o(S_s5_36_2), .c_out(C_s5_36_2));
logic S_s5_36_3, C_s5_36_3;
FA FA_s5_36_3(.A_i(C_s6_35_2), .B_i(C_s6_35_1), .c_in(C_s6_35_0), .S_o(S_s5_36_3), .c_out(C_s5_36_3));
logic S_s5_37_0, C_s5_37_0;
FA FA_s5_37_0(.A_i(S_s6_37_5), .B_i(S_s6_37_4), .c_in(S_s6_37_3), .S_o(S_s5_37_0), .c_out(C_s5_37_0));
logic S_s5_37_1, C_s5_37_1;
FA FA_s5_37_1(.A_i(S_s6_37_2), .B_i(S_s6_37_1), .c_in(S_s6_37_0), .S_o(S_s5_37_1), .c_out(C_s5_37_1));
logic S_s5_37_2, C_s5_37_2;
FA FA_s5_37_2(.A_i(C_s6_36_5), .B_i(C_s6_36_4), .c_in(C_s6_36_3), .S_o(S_s5_37_2), .c_out(C_s5_37_2));
logic S_s5_37_3, C_s5_37_3;
FA FA_s5_37_3(.A_i(C_s6_36_2), .B_i(C_s6_36_1), .c_in(C_s6_36_0), .S_o(S_s5_37_3), .c_out(C_s5_37_3));
logic S_s5_38_0, C_s5_38_0;
FA FA_s5_38_0(.A_i(S_s6_38_5), .B_i(S_s6_38_4), .c_in(S_s6_38_3), .S_o(S_s5_38_0), .c_out(C_s5_38_0));
logic S_s5_38_1, C_s5_38_1;
FA FA_s5_38_1(.A_i(S_s6_38_2), .B_i(S_s6_38_1), .c_in(S_s6_38_0), .S_o(S_s5_38_1), .c_out(C_s5_38_1));
logic S_s5_38_2, C_s5_38_2;
FA FA_s5_38_2(.A_i(C_s6_37_5), .B_i(C_s6_37_4), .c_in(C_s6_37_3), .S_o(S_s5_38_2), .c_out(C_s5_38_2));
logic S_s5_38_3, C_s5_38_3;
FA FA_s5_38_3(.A_i(C_s6_37_2), .B_i(C_s6_37_1), .c_in(C_s6_37_0), .S_o(S_s5_38_3), .c_out(C_s5_38_3));
logic S_s5_39_0, C_s5_39_0;
FA FA_s5_39_0(.A_i(S_s6_39_5), .B_i(S_s6_39_4), .c_in(S_s6_39_3), .S_o(S_s5_39_0), .c_out(C_s5_39_0));
logic S_s5_39_1, C_s5_39_1;
FA FA_s5_39_1(.A_i(S_s6_39_2), .B_i(S_s6_39_1), .c_in(S_s6_39_0), .S_o(S_s5_39_1), .c_out(C_s5_39_1));
logic S_s5_39_2, C_s5_39_2;
FA FA_s5_39_2(.A_i(C_s6_38_5), .B_i(C_s6_38_4), .c_in(C_s6_38_3), .S_o(S_s5_39_2), .c_out(C_s5_39_2));
logic S_s5_39_3, C_s5_39_3;
FA FA_s5_39_3(.A_i(C_s6_38_2), .B_i(C_s6_38_1), .c_in(C_s6_38_0), .S_o(S_s5_39_3), .c_out(C_s5_39_3));
logic S_s5_40_0, C_s5_40_0;
FA FA_s5_40_0(.A_i(S_s6_40_5), .B_i(S_s6_40_4), .c_in(S_s6_40_3), .S_o(S_s5_40_0), .c_out(C_s5_40_0));
logic S_s5_40_1, C_s5_40_1;
FA FA_s5_40_1(.A_i(S_s6_40_2), .B_i(S_s6_40_1), .c_in(S_s6_40_0), .S_o(S_s5_40_1), .c_out(C_s5_40_1));
logic S_s5_40_2, C_s5_40_2;
FA FA_s5_40_2(.A_i(C_s6_39_5), .B_i(C_s6_39_4), .c_in(C_s6_39_3), .S_o(S_s5_40_2), .c_out(C_s5_40_2));
logic S_s5_40_3, C_s5_40_3;
FA FA_s5_40_3(.A_i(C_s6_39_2), .B_i(C_s6_39_1), .c_in(C_s6_39_0), .S_o(S_s5_40_3), .c_out(C_s5_40_3));
logic S_s5_41_0, C_s5_41_0;
FA FA_s5_41_0(.A_i(S_s6_41_5), .B_i(S_s6_41_4), .c_in(S_s6_41_3), .S_o(S_s5_41_0), .c_out(C_s5_41_0));
logic S_s5_41_1, C_s5_41_1;
FA FA_s5_41_1(.A_i(S_s6_41_2), .B_i(S_s6_41_1), .c_in(S_s6_41_0), .S_o(S_s5_41_1), .c_out(C_s5_41_1));
logic S_s5_41_2, C_s5_41_2;
FA FA_s5_41_2(.A_i(C_s6_40_5), .B_i(C_s6_40_4), .c_in(C_s6_40_3), .S_o(S_s5_41_2), .c_out(C_s5_41_2));
logic S_s5_41_3, C_s5_41_3;
FA FA_s5_41_3(.A_i(C_s6_40_2), .B_i(C_s6_40_1), .c_in(C_s6_40_0), .S_o(S_s5_41_3), .c_out(C_s5_41_3));
logic S_s5_42_0, C_s5_42_0;
FA FA_s5_42_0(.A_i(S_s6_42_5), .B_i(S_s6_42_4), .c_in(S_s6_42_3), .S_o(S_s5_42_0), .c_out(C_s5_42_0));
logic S_s5_42_1, C_s5_42_1;
FA FA_s5_42_1(.A_i(S_s6_42_2), .B_i(S_s6_42_1), .c_in(S_s6_42_0), .S_o(S_s5_42_1), .c_out(C_s5_42_1));
logic S_s5_42_2, C_s5_42_2;
FA FA_s5_42_2(.A_i(C_s6_41_5), .B_i(C_s6_41_4), .c_in(C_s6_41_3), .S_o(S_s5_42_2), .c_out(C_s5_42_2));
logic S_s5_42_3, C_s5_42_3;
FA FA_s5_42_3(.A_i(C_s6_41_2), .B_i(C_s6_41_1), .c_in(C_s6_41_0), .S_o(S_s5_42_3), .c_out(C_s5_42_3));
logic S_s5_43_0, C_s5_43_0;
FA FA_s5_43_0(.A_i(S_s6_43_5), .B_i(S_s6_43_4), .c_in(S_s6_43_3), .S_o(S_s5_43_0), .c_out(C_s5_43_0));
logic S_s5_43_1, C_s5_43_1;
FA FA_s5_43_1(.A_i(S_s6_43_2), .B_i(S_s6_43_1), .c_in(S_s6_43_0), .S_o(S_s5_43_1), .c_out(C_s5_43_1));
logic S_s5_43_2, C_s5_43_2;
FA FA_s5_43_2(.A_i(C_s6_42_5), .B_i(C_s6_42_4), .c_in(C_s6_42_3), .S_o(S_s5_43_2), .c_out(C_s5_43_2));
logic S_s5_43_3, C_s5_43_3;
FA FA_s5_43_3(.A_i(C_s6_42_2), .B_i(C_s6_42_1), .c_in(C_s6_42_0), .S_o(S_s5_43_3), .c_out(C_s5_43_3));
logic S_s5_44_0, C_s5_44_0;
FA FA_s5_44_0(.A_i(S_s6_44_5), .B_i(S_s6_44_4), .c_in(S_s6_44_3), .S_o(S_s5_44_0), .c_out(C_s5_44_0));
logic S_s5_44_1, C_s5_44_1;
FA FA_s5_44_1(.A_i(S_s6_44_2), .B_i(S_s6_44_1), .c_in(S_s6_44_0), .S_o(S_s5_44_1), .c_out(C_s5_44_1));
logic S_s5_44_2, C_s5_44_2;
FA FA_s5_44_2(.A_i(C_s6_43_5), .B_i(C_s6_43_4), .c_in(C_s6_43_3), .S_o(S_s5_44_2), .c_out(C_s5_44_2));
logic S_s5_44_3, C_s5_44_3;
FA FA_s5_44_3(.A_i(C_s6_43_2), .B_i(C_s6_43_1), .c_in(C_s6_43_0), .S_o(S_s5_44_3), .c_out(C_s5_44_3));
logic S_s5_45_0, C_s5_45_0;
FA FA_s5_45_0(.A_i(S_s6_45_5), .B_i(S_s6_45_4), .c_in(S_s6_45_3), .S_o(S_s5_45_0), .c_out(C_s5_45_0));
logic S_s5_45_1, C_s5_45_1;
FA FA_s5_45_1(.A_i(S_s6_45_2), .B_i(S_s6_45_1), .c_in(S_s6_45_0), .S_o(S_s5_45_1), .c_out(C_s5_45_1));
logic S_s5_45_2, C_s5_45_2;
FA FA_s5_45_2(.A_i(C_s6_44_5), .B_i(C_s6_44_4), .c_in(C_s6_44_3), .S_o(S_s5_45_2), .c_out(C_s5_45_2));
logic S_s5_45_3, C_s5_45_3;
FA FA_s5_45_3(.A_i(C_s6_44_2), .B_i(C_s6_44_1), .c_in(C_s6_44_0), .S_o(S_s5_45_3), .c_out(C_s5_45_3));
logic S_s5_46_0, C_s5_46_0;
FA FA_s5_46_0(.A_i(S_s6_46_4), .B_i(S_s6_46_3), .c_in(S_s6_46_2), .S_o(S_s5_46_0), .c_out(C_s5_46_0));
logic S_s5_46_1, C_s5_46_1;
FA FA_s5_46_1(.A_i(S_s6_46_1), .B_i(S_s6_46_0), .c_in(C_s6_45_5), .S_o(S_s5_46_1), .c_out(C_s5_46_1));
logic S_s5_46_2, C_s5_46_2;
FA FA_s5_46_2(.A_i(C_s6_45_4), .B_i(C_s6_45_3), .c_in(C_s6_45_2), .S_o(S_s5_46_2), .c_out(C_s5_46_2));
logic S_s5_46_3, C_s5_46_3;
FA FA_s5_46_3(.A_i(C_s6_45_1), .B_i(C_s6_45_0), .c_in(comb[30][16]), .S_o(S_s5_46_3), .c_out(C_s5_46_3));
logic S_s5_47_0, C_s5_47_0;
FA FA_s5_47_0(.A_i(S_s6_47_3), .B_i(S_s6_47_2), .c_in(S_s6_47_1), .S_o(S_s5_47_0), .c_out(C_s5_47_0));
logic S_s5_47_1, C_s5_47_1;
FA FA_s5_47_1(.A_i(S_s6_47_0), .B_i(C_s6_46_4), .c_in(C_s6_46_3), .S_o(S_s5_47_1), .c_out(C_s5_47_1));
logic S_s5_47_2, C_s5_47_2;
FA FA_s5_47_2(.A_i(C_s6_46_2), .B_i(C_s6_46_1), .c_in(C_s6_46_0), .S_o(S_s5_47_2), .c_out(C_s5_47_2));
logic S_s5_47_3, C_s5_47_3;
FA FA_s5_47_3(.A_i(comb[28][19]), .B_i(comb[29][18]), .c_in(comb[30][17]), .S_o(S_s5_47_3), .c_out(C_s5_47_3));
logic S_s5_48_0, C_s5_48_0;
FA FA_s5_48_0(.A_i(S_s6_48_2), .B_i(S_s6_48_1), .c_in(S_s6_48_0), .S_o(S_s5_48_0), .c_out(C_s5_48_0));
logic S_s5_48_1, C_s5_48_1;
FA FA_s5_48_1(.A_i(C_s6_47_3), .B_i(C_s6_47_2), .c_in(C_s6_47_1), .S_o(S_s5_48_1), .c_out(C_s5_48_1));
logic S_s5_48_2, C_s5_48_2;
FA FA_s5_48_2(.A_i(C_s6_47_0), .B_i(comb[26][22]), .c_in(comb[27][21]), .S_o(S_s5_48_2), .c_out(C_s5_48_2));
logic S_s5_48_3, C_s5_48_3;
FA FA_s5_48_3(.A_i(comb[28][20]), .B_i(comb[29][19]), .c_in(comb[30][18]), .S_o(S_s5_48_3), .c_out(C_s5_48_3));
logic S_s5_49_0, C_s5_49_0;
FA FA_s5_49_0(.A_i(S_s6_49_1), .B_i(S_s6_49_0), .c_in(C_s6_48_2), .S_o(S_s5_49_0), .c_out(C_s5_49_0));
logic S_s5_49_1, C_s5_49_1;
FA FA_s5_49_1(.A_i(C_s6_48_1), .B_i(C_s6_48_0), .c_in(comb[24][25]), .S_o(S_s5_49_1), .c_out(C_s5_49_1));
logic S_s5_49_2, C_s5_49_2;
FA FA_s5_49_2(.A_i(comb[25][24]), .B_i(comb[26][23]), .c_in(comb[27][22]), .S_o(S_s5_49_2), .c_out(C_s5_49_2));
logic S_s5_49_3, C_s5_49_3;
FA FA_s5_49_3(.A_i(comb[28][21]), .B_i(comb[29][20]), .c_in(comb[30][19]), .S_o(S_s5_49_3), .c_out(C_s5_49_3));
logic S_s5_50_0, C_s5_50_0;
FA FA_s5_50_0(.A_i(S_s6_50_0), .B_i(C_s6_49_1), .c_in(C_s6_49_0), .S_o(S_s5_50_0), .c_out(C_s5_50_0));
logic S_s5_50_1, C_s5_50_1;
FA FA_s5_50_1(.A_i(comb[22][28]), .B_i(comb[23][27]), .c_in(comb[24][26]), .S_o(S_s5_50_1), .c_out(C_s5_50_1));
logic S_s5_50_2, C_s5_50_2;
FA FA_s5_50_2(.A_i(comb[25][25]), .B_i(comb[26][24]), .c_in(comb[27][23]), .S_o(S_s5_50_2), .c_out(C_s5_50_2));
logic S_s5_50_3, C_s5_50_3;
FA FA_s5_50_3(.A_i(comb[28][22]), .B_i(comb[29][21]), .c_in(comb[30][20]), .S_o(S_s5_50_3), .c_out(C_s5_50_3));
logic S_s5_51_0, C_s5_51_0;
FA FA_s5_51_0(.A_i(C_s6_50_0), .B_i(comb[20][31]), .c_in(comb[21][30]), .S_o(S_s5_51_0), .c_out(C_s5_51_0));
logic S_s5_51_1, C_s5_51_1;
FA FA_s5_51_1(.A_i(comb[22][29]), .B_i(comb[23][28]), .c_in(comb[24][27]), .S_o(S_s5_51_1), .c_out(C_s5_51_1));
logic S_s5_51_2, C_s5_51_2;
FA FA_s5_51_2(.A_i(comb[25][26]), .B_i(comb[26][25]), .c_in(comb[27][24]), .S_o(S_s5_51_2), .c_out(C_s5_51_2));
logic S_s5_51_3, C_s5_51_3;
FA FA_s5_51_3(.A_i(comb[28][23]), .B_i(comb[29][22]), .c_in(comb[30][21]), .S_o(S_s5_51_3), .c_out(C_s5_51_3));
logic S_s5_52_0, C_s5_52_0;
FA FA_s5_52_0(.A_i(comb[21][31]), .B_i(comb[22][30]), .c_in(comb[23][29]), .S_o(S_s5_52_0), .c_out(C_s5_52_0));
logic S_s5_52_1, C_s5_52_1;
FA FA_s5_52_1(.A_i(comb[24][28]), .B_i(comb[25][27]), .c_in(comb[26][26]), .S_o(S_s5_52_1), .c_out(C_s5_52_1));
logic S_s5_52_2, C_s5_52_2;
FA FA_s5_52_2(.A_i(comb[27][25]), .B_i(comb[28][24]), .c_in(comb[29][23]), .S_o(S_s5_52_2), .c_out(C_s5_52_2));
logic S_s5_53_0, C_s5_53_0;
FA FA_s5_53_0(.A_i(comb[22][31]), .B_i(comb[23][30]), .c_in(comb[24][29]), .S_o(S_s5_53_0), .c_out(C_s5_53_0));
logic S_s5_53_1, C_s5_53_1;
FA FA_s5_53_1(.A_i(comb[25][28]), .B_i(comb[26][27]), .c_in(comb[27][26]), .S_o(S_s5_53_1), .c_out(C_s5_53_1));
logic S_s5_54_0, C_s5_54_0;
FA FA_s5_54_0(.A_i(comb[23][31]), .B_i(comb[24][30]), .c_in(comb[25][29]), .S_o(S_s5_54_0), .c_out(C_s5_54_0));
// stage 5 end ======================================================================================================= 

// stage 4 begin ======================================================================================================= 
logic S_s4_6_0, C_s4_6_0;
HA HA_s4_60(.A_i(comb[0][6]), .B_i(comb[1][5]), .S_o(S_s4_6_0), .c_out(C_s4_6_0));
logic S_s4_7_0, C_s4_7_0;
FA FA_s4_7_0(.A_i(comb[0][7]), .B_i(comb[1][6]), .c_in(comb[2][5]), .S_o(S_s4_7_0), .c_out(C_s4_7_0));
logic S_s4_7_1, C_s4_7_1;
HA HA_s4_71(.A_i(comb[3][4]), .B_i(comb[4][3]), .S_o(S_s4_7_1), .c_out(C_s4_7_1));
logic S_s4_8_0, C_s4_8_0;
FA FA_s4_8_0(.A_i(comb[0][8]), .B_i(comb[1][7]), .c_in(comb[2][6]), .S_o(S_s4_8_0), .c_out(C_s4_8_0));
logic S_s4_8_1, C_s4_8_1;
FA FA_s4_8_1(.A_i(comb[3][5]), .B_i(comb[4][4]), .c_in(comb[5][3]), .S_o(S_s4_8_1), .c_out(C_s4_8_1));
logic S_s4_8_2, C_s4_8_2;
HA HA_s4_82(.A_i(comb[6][2]), .B_i(comb[7][1]), .S_o(S_s4_8_2), .c_out(C_s4_8_2));
logic S_s4_9_0, C_s4_9_0;
FA FA_s4_9_0(.A_i(S_s5_9_0), .B_i(comb[2][7]), .c_in(comb[3][6]), .S_o(S_s4_9_0), .c_out(C_s4_9_0));
logic S_s4_9_1, C_s4_9_1;
FA FA_s4_9_1(.A_i(comb[4][5]), .B_i(comb[5][4]), .c_in(comb[6][3]), .S_o(S_s4_9_1), .c_out(C_s4_9_1));
logic S_s4_9_2, C_s4_9_2;
FA FA_s4_9_2(.A_i(comb[7][2]), .B_i(comb[8][1]), .c_in(comb[9][0]), .S_o(S_s4_9_2), .c_out(C_s4_9_2));
logic S_s4_10_0, C_s4_10_0;
FA FA_s4_10_0(.A_i(S_s5_10_1), .B_i(S_s5_10_0), .c_in(C_s5_9_0), .S_o(S_s4_10_0), .c_out(C_s4_10_0));
logic S_s4_10_1, C_s4_10_1;
FA FA_s4_10_1(.A_i(comb[5][5]), .B_i(comb[6][4]), .c_in(comb[7][3]), .S_o(S_s4_10_1), .c_out(C_s4_10_1));
logic S_s4_10_2, C_s4_10_2;
FA FA_s4_10_2(.A_i(comb[8][2]), .B_i(comb[9][1]), .c_in(comb[10][0]), .S_o(S_s4_10_2), .c_out(C_s4_10_2));
logic S_s4_11_0, C_s4_11_0;
FA FA_s4_11_0(.A_i(S_s5_11_2), .B_i(S_s5_11_1), .c_in(S_s5_11_0), .S_o(S_s4_11_0), .c_out(C_s4_11_0));
logic S_s4_11_1, C_s4_11_1;
FA FA_s4_11_1(.A_i(C_s5_10_1), .B_i(C_s5_10_0), .c_in(comb[8][3]), .S_o(S_s4_11_1), .c_out(C_s4_11_1));
logic S_s4_11_2, C_s4_11_2;
FA FA_s4_11_2(.A_i(comb[9][2]), .B_i(comb[10][1]), .c_in(comb[11][0]), .S_o(S_s4_11_2), .c_out(C_s4_11_2));
logic S_s4_12_0, C_s4_12_0;
FA FA_s4_12_0(.A_i(S_s5_12_3), .B_i(S_s5_12_2), .c_in(S_s5_12_1), .S_o(S_s4_12_0), .c_out(C_s4_12_0));
logic S_s4_12_1, C_s4_12_1;
FA FA_s4_12_1(.A_i(S_s5_12_0), .B_i(C_s5_11_2), .c_in(C_s5_11_1), .S_o(S_s4_12_1), .c_out(C_s4_12_1));
logic S_s4_12_2, C_s4_12_2;
FA FA_s4_12_2(.A_i(C_s5_11_0), .B_i(comb[11][1]), .c_in(comb[12][0]), .S_o(S_s4_12_2), .c_out(C_s4_12_2));
logic S_s4_13_0, C_s4_13_0;
FA FA_s4_13_0(.A_i(S_s5_13_3), .B_i(S_s5_13_2), .c_in(S_s5_13_1), .S_o(S_s4_13_0), .c_out(C_s4_13_0));
logic S_s4_13_1, C_s4_13_1;
FA FA_s4_13_1(.A_i(S_s5_13_0), .B_i(C_s5_12_3), .c_in(C_s5_12_2), .S_o(S_s4_13_1), .c_out(C_s4_13_1));
logic S_s4_13_2, C_s4_13_2;
FA FA_s4_13_2(.A_i(C_s5_12_1), .B_i(C_s5_12_0), .c_in(comb[13][0]), .S_o(S_s4_13_2), .c_out(C_s4_13_2));
logic S_s4_14_0, C_s4_14_0;
FA FA_s4_14_0(.A_i(S_s5_14_3), .B_i(S_s5_14_2), .c_in(S_s5_14_1), .S_o(S_s4_14_0), .c_out(C_s4_14_0));
logic S_s4_14_1, C_s4_14_1;
FA FA_s4_14_1(.A_i(S_s5_14_0), .B_i(C_s5_13_3), .c_in(C_s5_13_2), .S_o(S_s4_14_1), .c_out(C_s4_14_1));
logic S_s4_14_2, C_s4_14_2;
FA FA_s4_14_2(.A_i(C_s5_13_1), .B_i(C_s5_13_0), .c_in(comb[14][0]), .S_o(S_s4_14_2), .c_out(C_s4_14_2));
logic S_s4_15_0, C_s4_15_0;
FA FA_s4_15_0(.A_i(S_s5_15_3), .B_i(S_s5_15_2), .c_in(S_s5_15_1), .S_o(S_s4_15_0), .c_out(C_s4_15_0));
logic S_s4_15_1, C_s4_15_1;
FA FA_s4_15_1(.A_i(S_s5_15_0), .B_i(C_s5_14_3), .c_in(C_s5_14_2), .S_o(S_s4_15_1), .c_out(C_s4_15_1));
logic S_s4_15_2, C_s4_15_2;
FA FA_s4_15_2(.A_i(C_s5_14_1), .B_i(C_s5_14_0), .c_in(comb[15][0]), .S_o(S_s4_15_2), .c_out(C_s4_15_2));
logic S_s4_16_0, C_s4_16_0;
FA FA_s4_16_0(.A_i(S_s5_16_3), .B_i(S_s5_16_2), .c_in(S_s5_16_1), .S_o(S_s4_16_0), .c_out(C_s4_16_0));
logic S_s4_16_1, C_s4_16_1;
FA FA_s4_16_1(.A_i(S_s5_16_0), .B_i(C_s5_15_3), .c_in(C_s5_15_2), .S_o(S_s4_16_1), .c_out(C_s4_16_1));
logic S_s4_16_2, C_s4_16_2;
FA FA_s4_16_2(.A_i(C_s5_15_1), .B_i(C_s5_15_0), .c_in(comb[16][0]), .S_o(S_s4_16_2), .c_out(C_s4_16_2));
logic S_s4_17_0, C_s4_17_0;
FA FA_s4_17_0(.A_i(S_s5_17_3), .B_i(S_s5_17_2), .c_in(S_s5_17_1), .S_o(S_s4_17_0), .c_out(C_s4_17_0));
logic S_s4_17_1, C_s4_17_1;
FA FA_s4_17_1(.A_i(S_s5_17_0), .B_i(C_s5_16_3), .c_in(C_s5_16_2), .S_o(S_s4_17_1), .c_out(C_s4_17_1));
logic S_s4_17_2, C_s4_17_2;
FA FA_s4_17_2(.A_i(C_s5_16_1), .B_i(C_s5_16_0), .c_in(comb[17][0]), .S_o(S_s4_17_2), .c_out(C_s4_17_2));
logic S_s4_18_0, C_s4_18_0;
FA FA_s4_18_0(.A_i(S_s5_18_3), .B_i(S_s5_18_2), .c_in(S_s5_18_1), .S_o(S_s4_18_0), .c_out(C_s4_18_0));
logic S_s4_18_1, C_s4_18_1;
FA FA_s4_18_1(.A_i(S_s5_18_0), .B_i(C_s5_17_3), .c_in(C_s5_17_2), .S_o(S_s4_18_1), .c_out(C_s4_18_1));
logic S_s4_18_2, C_s4_18_2;
FA FA_s4_18_2(.A_i(C_s5_17_1), .B_i(C_s5_17_0), .c_in(comb[18][0]), .S_o(S_s4_18_2), .c_out(C_s4_18_2));
logic S_s4_19_0, C_s4_19_0;
FA FA_s4_19_0(.A_i(S_s5_19_3), .B_i(S_s5_19_2), .c_in(S_s5_19_1), .S_o(S_s4_19_0), .c_out(C_s4_19_0));
logic S_s4_19_1, C_s4_19_1;
FA FA_s4_19_1(.A_i(S_s5_19_0), .B_i(C_s5_18_3), .c_in(C_s5_18_2), .S_o(S_s4_19_1), .c_out(C_s4_19_1));
logic S_s4_19_2, C_s4_19_2;
FA FA_s4_19_2(.A_i(C_s5_18_1), .B_i(C_s5_18_0), .c_in(comb[19][0]), .S_o(S_s4_19_2), .c_out(C_s4_19_2));
logic S_s4_20_0, C_s4_20_0;
FA FA_s4_20_0(.A_i(S_s5_20_3), .B_i(S_s5_20_2), .c_in(S_s5_20_1), .S_o(S_s4_20_0), .c_out(C_s4_20_0));
logic S_s4_20_1, C_s4_20_1;
FA FA_s4_20_1(.A_i(S_s5_20_0), .B_i(C_s5_19_3), .c_in(C_s5_19_2), .S_o(S_s4_20_1), .c_out(C_s4_20_1));
logic S_s4_20_2, C_s4_20_2;
FA FA_s4_20_2(.A_i(C_s5_19_1), .B_i(C_s5_19_0), .c_in(comb[20][0]), .S_o(S_s4_20_2), .c_out(C_s4_20_2));
logic S_s4_21_0, C_s4_21_0;
FA FA_s4_21_0(.A_i(S_s5_21_3), .B_i(S_s5_21_2), .c_in(S_s5_21_1), .S_o(S_s4_21_0), .c_out(C_s4_21_0));
logic S_s4_21_1, C_s4_21_1;
FA FA_s4_21_1(.A_i(S_s5_21_0), .B_i(C_s5_20_3), .c_in(C_s5_20_2), .S_o(S_s4_21_1), .c_out(C_s4_21_1));
logic S_s4_21_2, C_s4_21_2;
FA FA_s4_21_2(.A_i(C_s5_20_1), .B_i(C_s5_20_0), .c_in(comb[21][0]), .S_o(S_s4_21_2), .c_out(C_s4_21_2));
logic S_s4_22_0, C_s4_22_0;
FA FA_s4_22_0(.A_i(S_s5_22_3), .B_i(S_s5_22_2), .c_in(S_s5_22_1), .S_o(S_s4_22_0), .c_out(C_s4_22_0));
logic S_s4_22_1, C_s4_22_1;
FA FA_s4_22_1(.A_i(S_s5_22_0), .B_i(C_s5_21_3), .c_in(C_s5_21_2), .S_o(S_s4_22_1), .c_out(C_s4_22_1));
logic S_s4_22_2, C_s4_22_2;
FA FA_s4_22_2(.A_i(C_s5_21_1), .B_i(C_s5_21_0), .c_in(comb[22][0]), .S_o(S_s4_22_2), .c_out(C_s4_22_2));
logic S_s4_23_0, C_s4_23_0;
FA FA_s4_23_0(.A_i(S_s5_23_3), .B_i(S_s5_23_2), .c_in(S_s5_23_1), .S_o(S_s4_23_0), .c_out(C_s4_23_0));
logic S_s4_23_1, C_s4_23_1;
FA FA_s4_23_1(.A_i(S_s5_23_0), .B_i(C_s5_22_3), .c_in(C_s5_22_2), .S_o(S_s4_23_1), .c_out(C_s4_23_1));
logic S_s4_23_2, C_s4_23_2;
FA FA_s4_23_2(.A_i(C_s5_22_1), .B_i(C_s5_22_0), .c_in(comb[23][0]), .S_o(S_s4_23_2), .c_out(C_s4_23_2));
logic S_s4_24_0, C_s4_24_0;
FA FA_s4_24_0(.A_i(S_s5_24_3), .B_i(S_s5_24_2), .c_in(S_s5_24_1), .S_o(S_s4_24_0), .c_out(C_s4_24_0));
logic S_s4_24_1, C_s4_24_1;
FA FA_s4_24_1(.A_i(S_s5_24_0), .B_i(C_s5_23_3), .c_in(C_s5_23_2), .S_o(S_s4_24_1), .c_out(C_s4_24_1));
logic S_s4_24_2, C_s4_24_2;
FA FA_s4_24_2(.A_i(C_s5_23_1), .B_i(C_s5_23_0), .c_in(comb[24][0]), .S_o(S_s4_24_2), .c_out(C_s4_24_2));
logic S_s4_25_0, C_s4_25_0;
FA FA_s4_25_0(.A_i(S_s5_25_3), .B_i(S_s5_25_2), .c_in(S_s5_25_1), .S_o(S_s4_25_0), .c_out(C_s4_25_0));
logic S_s4_25_1, C_s4_25_1;
FA FA_s4_25_1(.A_i(S_s5_25_0), .B_i(C_s5_24_3), .c_in(C_s5_24_2), .S_o(S_s4_25_1), .c_out(C_s4_25_1));
logic S_s4_25_2, C_s4_25_2;
FA FA_s4_25_2(.A_i(C_s5_24_1), .B_i(C_s5_24_0), .c_in(comb[25][0]), .S_o(S_s4_25_2), .c_out(C_s4_25_2));
logic S_s4_26_0, C_s4_26_0;
FA FA_s4_26_0(.A_i(S_s5_26_3), .B_i(S_s5_26_2), .c_in(S_s5_26_1), .S_o(S_s4_26_0), .c_out(C_s4_26_0));
logic S_s4_26_1, C_s4_26_1;
FA FA_s4_26_1(.A_i(S_s5_26_0), .B_i(C_s5_25_3), .c_in(C_s5_25_2), .S_o(S_s4_26_1), .c_out(C_s4_26_1));
logic S_s4_26_2, C_s4_26_2;
FA FA_s4_26_2(.A_i(C_s5_25_1), .B_i(C_s5_25_0), .c_in(comb[26][0]), .S_o(S_s4_26_2), .c_out(C_s4_26_2));
logic S_s4_27_0, C_s4_27_0;
FA FA_s4_27_0(.A_i(S_s5_27_3), .B_i(S_s5_27_2), .c_in(S_s5_27_1), .S_o(S_s4_27_0), .c_out(C_s4_27_0));
logic S_s4_27_1, C_s4_27_1;
FA FA_s4_27_1(.A_i(S_s5_27_0), .B_i(C_s5_26_3), .c_in(C_s5_26_2), .S_o(S_s4_27_1), .c_out(C_s4_27_1));
logic S_s4_27_2, C_s4_27_2;
FA FA_s4_27_2(.A_i(C_s5_26_1), .B_i(C_s5_26_0), .c_in(comb[27][0]), .S_o(S_s4_27_2), .c_out(C_s4_27_2));
logic S_s4_28_0, C_s4_28_0;
FA FA_s4_28_0(.A_i(S_s5_28_3), .B_i(S_s5_28_2), .c_in(S_s5_28_1), .S_o(S_s4_28_0), .c_out(C_s4_28_0));
logic S_s4_28_1, C_s4_28_1;
FA FA_s4_28_1(.A_i(S_s5_28_0), .B_i(C_s5_27_3), .c_in(C_s5_27_2), .S_o(S_s4_28_1), .c_out(C_s4_28_1));
logic S_s4_28_2, C_s4_28_2;
FA FA_s4_28_2(.A_i(C_s5_27_1), .B_i(C_s5_27_0), .c_in(comb[28][0]), .S_o(S_s4_28_2), .c_out(C_s4_28_2));
logic S_s4_29_0, C_s4_29_0;
FA FA_s4_29_0(.A_i(S_s5_29_3), .B_i(S_s5_29_2), .c_in(S_s5_29_1), .S_o(S_s4_29_0), .c_out(C_s4_29_0));
logic S_s4_29_1, C_s4_29_1;
FA FA_s4_29_1(.A_i(S_s5_29_0), .B_i(C_s5_28_3), .c_in(C_s5_28_2), .S_o(S_s4_29_1), .c_out(C_s4_29_1));
logic S_s4_29_2, C_s4_29_2;
FA FA_s4_29_2(.A_i(C_s5_28_1), .B_i(C_s5_28_0), .c_in(comb[29][0]), .S_o(S_s4_29_2), .c_out(C_s4_29_2));
logic S_s4_30_0, C_s4_30_0;
FA FA_s4_30_0(.A_i(S_s5_30_3), .B_i(S_s5_30_2), .c_in(S_s5_30_1), .S_o(S_s4_30_0), .c_out(C_s4_30_0));
logic S_s4_30_1, C_s4_30_1;
FA FA_s4_30_1(.A_i(S_s5_30_0), .B_i(C_s5_29_3), .c_in(C_s5_29_2), .S_o(S_s4_30_1), .c_out(C_s4_30_1));
logic S_s4_30_2, C_s4_30_2;
FA FA_s4_30_2(.A_i(C_s5_29_1), .B_i(C_s5_29_0), .c_in(comb[30][0]), .S_o(S_s4_30_2), .c_out(C_s4_30_2));
logic S_s4_31_0, C_s4_31_0;
FA FA_s4_31_0(.A_i(S_s5_31_3), .B_i(S_s5_31_2), .c_in(S_s5_31_1), .S_o(S_s4_31_0), .c_out(C_s4_31_0));
logic S_s4_31_1, C_s4_31_1;
FA FA_s4_31_1(.A_i(S_s5_31_0), .B_i(C_s5_30_3), .c_in(C_s5_30_2), .S_o(S_s4_31_1), .c_out(C_s4_31_1));
logic S_s4_31_2, C_s4_31_2;
FA FA_s4_31_2(.A_i(C_s5_30_1), .B_i(C_s5_30_0), .c_in(comb[31][0]), .S_o(S_s4_31_2), .c_out(C_s4_31_2));
logic S_s4_32_0, C_s4_32_0;
FA FA_s4_32_0(.A_i(S_s5_32_3), .B_i(S_s5_32_2), .c_in(S_s5_32_1), .S_o(S_s4_32_0), .c_out(C_s4_32_0));
logic S_s4_32_1, C_s4_32_1;
FA FA_s4_32_1(.A_i(S_s5_32_0), .B_i(C_s5_31_3), .c_in(C_s5_31_2), .S_o(S_s4_32_1), .c_out(C_s4_32_1));
logic S_s4_32_2, C_s4_32_2;
FA FA_s4_32_2(.A_i(C_s5_31_1), .B_i(C_s5_31_0), .c_in(comb[31][1]), .S_o(S_s4_32_2), .c_out(C_s4_32_2));
logic S_s4_33_0, C_s4_33_0;
FA FA_s4_33_0(.A_i(S_s5_33_3), .B_i(S_s5_33_2), .c_in(S_s5_33_1), .S_o(S_s4_33_0), .c_out(C_s4_33_0));
logic S_s4_33_1, C_s4_33_1;
FA FA_s4_33_1(.A_i(S_s5_33_0), .B_i(C_s5_32_3), .c_in(C_s5_32_2), .S_o(S_s4_33_1), .c_out(C_s4_33_1));
logic S_s4_33_2, C_s4_33_2;
FA FA_s4_33_2(.A_i(C_s5_32_1), .B_i(C_s5_32_0), .c_in(comb[31][2]), .S_o(S_s4_33_2), .c_out(C_s4_33_2));
logic S_s4_34_0, C_s4_34_0;
FA FA_s4_34_0(.A_i(S_s5_34_3), .B_i(S_s5_34_2), .c_in(S_s5_34_1), .S_o(S_s4_34_0), .c_out(C_s4_34_0));
logic S_s4_34_1, C_s4_34_1;
FA FA_s4_34_1(.A_i(S_s5_34_0), .B_i(C_s5_33_3), .c_in(C_s5_33_2), .S_o(S_s4_34_1), .c_out(C_s4_34_1));
logic S_s4_34_2, C_s4_34_2;
FA FA_s4_34_2(.A_i(C_s5_33_1), .B_i(C_s5_33_0), .c_in(comb[31][3]), .S_o(S_s4_34_2), .c_out(C_s4_34_2));
logic S_s4_35_0, C_s4_35_0;
FA FA_s4_35_0(.A_i(S_s5_35_3), .B_i(S_s5_35_2), .c_in(S_s5_35_1), .S_o(S_s4_35_0), .c_out(C_s4_35_0));
logic S_s4_35_1, C_s4_35_1;
FA FA_s4_35_1(.A_i(S_s5_35_0), .B_i(C_s5_34_3), .c_in(C_s5_34_2), .S_o(S_s4_35_1), .c_out(C_s4_35_1));
logic S_s4_35_2, C_s4_35_2;
FA FA_s4_35_2(.A_i(C_s5_34_1), .B_i(C_s5_34_0), .c_in(comb[31][4]), .S_o(S_s4_35_2), .c_out(C_s4_35_2));
logic S_s4_36_0, C_s4_36_0;
FA FA_s4_36_0(.A_i(S_s5_36_3), .B_i(S_s5_36_2), .c_in(S_s5_36_1), .S_o(S_s4_36_0), .c_out(C_s4_36_0));
logic S_s4_36_1, C_s4_36_1;
FA FA_s4_36_1(.A_i(S_s5_36_0), .B_i(C_s5_35_3), .c_in(C_s5_35_2), .S_o(S_s4_36_1), .c_out(C_s4_36_1));
logic S_s4_36_2, C_s4_36_2;
FA FA_s4_36_2(.A_i(C_s5_35_1), .B_i(C_s5_35_0), .c_in(comb[31][5]), .S_o(S_s4_36_2), .c_out(C_s4_36_2));
logic S_s4_37_0, C_s4_37_0;
FA FA_s4_37_0(.A_i(S_s5_37_3), .B_i(S_s5_37_2), .c_in(S_s5_37_1), .S_o(S_s4_37_0), .c_out(C_s4_37_0));
logic S_s4_37_1, C_s4_37_1;
FA FA_s4_37_1(.A_i(S_s5_37_0), .B_i(C_s5_36_3), .c_in(C_s5_36_2), .S_o(S_s4_37_1), .c_out(C_s4_37_1));
logic S_s4_37_2, C_s4_37_2;
FA FA_s4_37_2(.A_i(C_s5_36_1), .B_i(C_s5_36_0), .c_in(comb[31][6]), .S_o(S_s4_37_2), .c_out(C_s4_37_2));
logic S_s4_38_0, C_s4_38_0;
FA FA_s4_38_0(.A_i(S_s5_38_3), .B_i(S_s5_38_2), .c_in(S_s5_38_1), .S_o(S_s4_38_0), .c_out(C_s4_38_0));
logic S_s4_38_1, C_s4_38_1;
FA FA_s4_38_1(.A_i(S_s5_38_0), .B_i(C_s5_37_3), .c_in(C_s5_37_2), .S_o(S_s4_38_1), .c_out(C_s4_38_1));
logic S_s4_38_2, C_s4_38_2;
FA FA_s4_38_2(.A_i(C_s5_37_1), .B_i(C_s5_37_0), .c_in(comb[31][7]), .S_o(S_s4_38_2), .c_out(C_s4_38_2));
logic S_s4_39_0, C_s4_39_0;
FA FA_s4_39_0(.A_i(S_s5_39_3), .B_i(S_s5_39_2), .c_in(S_s5_39_1), .S_o(S_s4_39_0), .c_out(C_s4_39_0));
logic S_s4_39_1, C_s4_39_1;
FA FA_s4_39_1(.A_i(S_s5_39_0), .B_i(C_s5_38_3), .c_in(C_s5_38_2), .S_o(S_s4_39_1), .c_out(C_s4_39_1));
logic S_s4_39_2, C_s4_39_2;
FA FA_s4_39_2(.A_i(C_s5_38_1), .B_i(C_s5_38_0), .c_in(comb[31][8]), .S_o(S_s4_39_2), .c_out(C_s4_39_2));
logic S_s4_40_0, C_s4_40_0;
FA FA_s4_40_0(.A_i(S_s5_40_3), .B_i(S_s5_40_2), .c_in(S_s5_40_1), .S_o(S_s4_40_0), .c_out(C_s4_40_0));
logic S_s4_40_1, C_s4_40_1;
FA FA_s4_40_1(.A_i(S_s5_40_0), .B_i(C_s5_39_3), .c_in(C_s5_39_2), .S_o(S_s4_40_1), .c_out(C_s4_40_1));
logic S_s4_40_2, C_s4_40_2;
FA FA_s4_40_2(.A_i(C_s5_39_1), .B_i(C_s5_39_0), .c_in(comb[31][9]), .S_o(S_s4_40_2), .c_out(C_s4_40_2));
logic S_s4_41_0, C_s4_41_0;
FA FA_s4_41_0(.A_i(S_s5_41_3), .B_i(S_s5_41_2), .c_in(S_s5_41_1), .S_o(S_s4_41_0), .c_out(C_s4_41_0));
logic S_s4_41_1, C_s4_41_1;
FA FA_s4_41_1(.A_i(S_s5_41_0), .B_i(C_s5_40_3), .c_in(C_s5_40_2), .S_o(S_s4_41_1), .c_out(C_s4_41_1));
logic S_s4_41_2, C_s4_41_2;
FA FA_s4_41_2(.A_i(C_s5_40_1), .B_i(C_s5_40_0), .c_in(comb[31][10]), .S_o(S_s4_41_2), .c_out(C_s4_41_2));
logic S_s4_42_0, C_s4_42_0;
FA FA_s4_42_0(.A_i(S_s5_42_3), .B_i(S_s5_42_2), .c_in(S_s5_42_1), .S_o(S_s4_42_0), .c_out(C_s4_42_0));
logic S_s4_42_1, C_s4_42_1;
FA FA_s4_42_1(.A_i(S_s5_42_0), .B_i(C_s5_41_3), .c_in(C_s5_41_2), .S_o(S_s4_42_1), .c_out(C_s4_42_1));
logic S_s4_42_2, C_s4_42_2;
FA FA_s4_42_2(.A_i(C_s5_41_1), .B_i(C_s5_41_0), .c_in(comb[31][11]), .S_o(S_s4_42_2), .c_out(C_s4_42_2));
logic S_s4_43_0, C_s4_43_0;
FA FA_s4_43_0(.A_i(S_s5_43_3), .B_i(S_s5_43_2), .c_in(S_s5_43_1), .S_o(S_s4_43_0), .c_out(C_s4_43_0));
logic S_s4_43_1, C_s4_43_1;
FA FA_s4_43_1(.A_i(S_s5_43_0), .B_i(C_s5_42_3), .c_in(C_s5_42_2), .S_o(S_s4_43_1), .c_out(C_s4_43_1));
logic S_s4_43_2, C_s4_43_2;
FA FA_s4_43_2(.A_i(C_s5_42_1), .B_i(C_s5_42_0), .c_in(comb[31][12]), .S_o(S_s4_43_2), .c_out(C_s4_43_2));
logic S_s4_44_0, C_s4_44_0;
FA FA_s4_44_0(.A_i(S_s5_44_3), .B_i(S_s5_44_2), .c_in(S_s5_44_1), .S_o(S_s4_44_0), .c_out(C_s4_44_0));
logic S_s4_44_1, C_s4_44_1;
FA FA_s4_44_1(.A_i(S_s5_44_0), .B_i(C_s5_43_3), .c_in(C_s5_43_2), .S_o(S_s4_44_1), .c_out(C_s4_44_1));
logic S_s4_44_2, C_s4_44_2;
FA FA_s4_44_2(.A_i(C_s5_43_1), .B_i(C_s5_43_0), .c_in(comb[31][13]), .S_o(S_s4_44_2), .c_out(C_s4_44_2));
logic S_s4_45_0, C_s4_45_0;
FA FA_s4_45_0(.A_i(S_s5_45_3), .B_i(S_s5_45_2), .c_in(S_s5_45_1), .S_o(S_s4_45_0), .c_out(C_s4_45_0));
logic S_s4_45_1, C_s4_45_1;
FA FA_s4_45_1(.A_i(S_s5_45_0), .B_i(C_s5_44_3), .c_in(C_s5_44_2), .S_o(S_s4_45_1), .c_out(C_s4_45_1));
logic S_s4_45_2, C_s4_45_2;
FA FA_s4_45_2(.A_i(C_s5_44_1), .B_i(C_s5_44_0), .c_in(comb[31][14]), .S_o(S_s4_45_2), .c_out(C_s4_45_2));
logic S_s4_46_0, C_s4_46_0;
FA FA_s4_46_0(.A_i(S_s5_46_3), .B_i(S_s5_46_2), .c_in(S_s5_46_1), .S_o(S_s4_46_0), .c_out(C_s4_46_0));
logic S_s4_46_1, C_s4_46_1;
FA FA_s4_46_1(.A_i(S_s5_46_0), .B_i(C_s5_45_3), .c_in(C_s5_45_2), .S_o(S_s4_46_1), .c_out(C_s4_46_1));
logic S_s4_46_2, C_s4_46_2;
FA FA_s4_46_2(.A_i(C_s5_45_1), .B_i(C_s5_45_0), .c_in(comb[31][15]), .S_o(S_s4_46_2), .c_out(C_s4_46_2));
logic S_s4_47_0, C_s4_47_0;
FA FA_s4_47_0(.A_i(S_s5_47_3), .B_i(S_s5_47_2), .c_in(S_s5_47_1), .S_o(S_s4_47_0), .c_out(C_s4_47_0));
logic S_s4_47_1, C_s4_47_1;
FA FA_s4_47_1(.A_i(S_s5_47_0), .B_i(C_s5_46_3), .c_in(C_s5_46_2), .S_o(S_s4_47_1), .c_out(C_s4_47_1));
logic S_s4_47_2, C_s4_47_2;
FA FA_s4_47_2(.A_i(C_s5_46_1), .B_i(C_s5_46_0), .c_in(comb[31][16]), .S_o(S_s4_47_2), .c_out(C_s4_47_2));
logic S_s4_48_0, C_s4_48_0;
FA FA_s4_48_0(.A_i(S_s5_48_3), .B_i(S_s5_48_2), .c_in(S_s5_48_1), .S_o(S_s4_48_0), .c_out(C_s4_48_0));
logic S_s4_48_1, C_s4_48_1;
FA FA_s4_48_1(.A_i(S_s5_48_0), .B_i(C_s5_47_3), .c_in(C_s5_47_2), .S_o(S_s4_48_1), .c_out(C_s4_48_1));
logic S_s4_48_2, C_s4_48_2;
FA FA_s4_48_2(.A_i(C_s5_47_1), .B_i(C_s5_47_0), .c_in(comb[31][17]), .S_o(S_s4_48_2), .c_out(C_s4_48_2));
logic S_s4_49_0, C_s4_49_0;
FA FA_s4_49_0(.A_i(S_s5_49_3), .B_i(S_s5_49_2), .c_in(S_s5_49_1), .S_o(S_s4_49_0), .c_out(C_s4_49_0));
logic S_s4_49_1, C_s4_49_1;
FA FA_s4_49_1(.A_i(S_s5_49_0), .B_i(C_s5_48_3), .c_in(C_s5_48_2), .S_o(S_s4_49_1), .c_out(C_s4_49_1));
logic S_s4_49_2, C_s4_49_2;
FA FA_s4_49_2(.A_i(C_s5_48_1), .B_i(C_s5_48_0), .c_in(comb[31][18]), .S_o(S_s4_49_2), .c_out(C_s4_49_2));
logic S_s4_50_0, C_s4_50_0;
FA FA_s4_50_0(.A_i(S_s5_50_3), .B_i(S_s5_50_2), .c_in(S_s5_50_1), .S_o(S_s4_50_0), .c_out(C_s4_50_0));
logic S_s4_50_1, C_s4_50_1;
FA FA_s4_50_1(.A_i(S_s5_50_0), .B_i(C_s5_49_3), .c_in(C_s5_49_2), .S_o(S_s4_50_1), .c_out(C_s4_50_1));
logic S_s4_50_2, C_s4_50_2;
FA FA_s4_50_2(.A_i(C_s5_49_1), .B_i(C_s5_49_0), .c_in(comb[31][19]), .S_o(S_s4_50_2), .c_out(C_s4_50_2));
logic S_s4_51_0, C_s4_51_0;
FA FA_s4_51_0(.A_i(S_s5_51_3), .B_i(S_s5_51_2), .c_in(S_s5_51_1), .S_o(S_s4_51_0), .c_out(C_s4_51_0));
logic S_s4_51_1, C_s4_51_1;
FA FA_s4_51_1(.A_i(S_s5_51_0), .B_i(C_s5_50_3), .c_in(C_s5_50_2), .S_o(S_s4_51_1), .c_out(C_s4_51_1));
logic S_s4_51_2, C_s4_51_2;
FA FA_s4_51_2(.A_i(C_s5_50_1), .B_i(C_s5_50_0), .c_in(comb[31][20]), .S_o(S_s4_51_2), .c_out(C_s4_51_2));
logic S_s4_52_0, C_s4_52_0;
FA FA_s4_52_0(.A_i(S_s5_52_2), .B_i(S_s5_52_1), .c_in(S_s5_52_0), .S_o(S_s4_52_0), .c_out(C_s4_52_0));
logic S_s4_52_1, C_s4_52_1;
FA FA_s4_52_1(.A_i(C_s5_51_3), .B_i(C_s5_51_2), .c_in(C_s5_51_1), .S_o(S_s4_52_1), .c_out(C_s4_52_1));
logic S_s4_52_2, C_s4_52_2;
FA FA_s4_52_2(.A_i(C_s5_51_0), .B_i(comb[30][22]), .c_in(comb[31][21]), .S_o(S_s4_52_2), .c_out(C_s4_52_2));
logic S_s4_53_0, C_s4_53_0;
FA FA_s4_53_0(.A_i(S_s5_53_1), .B_i(S_s5_53_0), .c_in(C_s5_52_2), .S_o(S_s4_53_0), .c_out(C_s4_53_0));
logic S_s4_53_1, C_s4_53_1;
FA FA_s4_53_1(.A_i(C_s5_52_1), .B_i(C_s5_52_0), .c_in(comb[28][25]), .S_o(S_s4_53_1), .c_out(C_s4_53_1));
logic S_s4_53_2, C_s4_53_2;
FA FA_s4_53_2(.A_i(comb[29][24]), .B_i(comb[30][23]), .c_in(comb[31][22]), .S_o(S_s4_53_2), .c_out(C_s4_53_2));
logic S_s4_54_0, C_s4_54_0;
FA FA_s4_54_0(.A_i(S_s5_54_0), .B_i(C_s5_53_1), .c_in(C_s5_53_0), .S_o(S_s4_54_0), .c_out(C_s4_54_0));
logic S_s4_54_1, C_s4_54_1;
FA FA_s4_54_1(.A_i(comb[26][28]), .B_i(comb[27][27]), .c_in(comb[28][26]), .S_o(S_s4_54_1), .c_out(C_s4_54_1));
logic S_s4_54_2, C_s4_54_2;
FA FA_s4_54_2(.A_i(comb[29][25]), .B_i(comb[30][24]), .c_in(comb[31][23]), .S_o(S_s4_54_2), .c_out(C_s4_54_2));
logic S_s4_55_0, C_s4_55_0;
FA FA_s4_55_0(.A_i(C_s5_54_0), .B_i(comb[24][31]), .c_in(comb[25][30]), .S_o(S_s4_55_0), .c_out(C_s4_55_0));
logic S_s4_55_1, C_s4_55_1;
FA FA_s4_55_1(.A_i(comb[26][29]), .B_i(comb[27][28]), .c_in(comb[28][27]), .S_o(S_s4_55_1), .c_out(C_s4_55_1));
logic S_s4_55_2, C_s4_55_2;
FA FA_s4_55_2(.A_i(comb[29][26]), .B_i(comb[30][25]), .c_in(comb[31][24]), .S_o(S_s4_55_2), .c_out(C_s4_55_2));
logic S_s4_56_0, C_s4_56_0;
FA FA_s4_56_0(.A_i(comb[25][31]), .B_i(comb[26][30]), .c_in(comb[27][29]), .S_o(S_s4_56_0), .c_out(C_s4_56_0));
logic S_s4_56_1, C_s4_56_1;
FA FA_s4_56_1(.A_i(comb[28][28]), .B_i(comb[29][27]), .c_in(comb[30][26]), .S_o(S_s4_56_1), .c_out(C_s4_56_1));
logic S_s4_57_0, C_s4_57_0;
FA FA_s4_57_0(.A_i(comb[26][31]), .B_i(comb[27][30]), .c_in(comb[28][29]), .S_o(S_s4_57_0), .c_out(C_s4_57_0));
// stage 4 end ======================================================================================================= 

// stage 3 begin ======================================================================================================= 
logic S_s3_4_0, C_s3_4_0;
HA HA_s3_40(.A_i(comb[0][4]), .B_i(comb[1][3]), .S_o(S_s3_4_0), .c_out(C_s3_4_0));
logic S_s3_5_0, C_s3_5_0;
FA FA_s3_5_0(.A_i(comb[0][5]), .B_i(comb[1][4]), .c_in(comb[2][3]), .S_o(S_s3_5_0), .c_out(C_s3_5_0));
logic S_s3_5_1, C_s3_5_1;
HA HA_s3_51(.A_i(comb[3][2]), .B_i(comb[4][1]), .S_o(S_s3_5_1), .c_out(C_s3_5_1));
logic S_s3_6_0, C_s3_6_0;
FA FA_s3_6_0(.A_i(S_s4_6_0), .B_i(comb[2][4]), .c_in(comb[3][3]), .S_o(S_s3_6_0), .c_out(C_s3_6_0));
logic S_s3_6_1, C_s3_6_1;
FA FA_s3_6_1(.A_i(comb[4][2]), .B_i(comb[5][1]), .c_in(comb[6][0]), .S_o(S_s3_6_1), .c_out(C_s3_6_1));
logic S_s3_7_0, C_s3_7_0;
FA FA_s3_7_0(.A_i(S_s4_7_1), .B_i(S_s4_7_0), .c_in(C_s4_6_0), .S_o(S_s3_7_0), .c_out(C_s3_7_0));
logic S_s3_7_1, C_s3_7_1;
FA FA_s3_7_1(.A_i(comb[5][2]), .B_i(comb[6][1]), .c_in(comb[7][0]), .S_o(S_s3_7_1), .c_out(C_s3_7_1));
logic S_s3_8_0, C_s3_8_0;
FA FA_s3_8_0(.A_i(S_s4_8_2), .B_i(S_s4_8_1), .c_in(S_s4_8_0), .S_o(S_s3_8_0), .c_out(C_s3_8_0));
logic S_s3_8_1, C_s3_8_1;
FA FA_s3_8_1(.A_i(C_s4_7_1), .B_i(C_s4_7_0), .c_in(comb[8][0]), .S_o(S_s3_8_1), .c_out(C_s3_8_1));
logic S_s3_9_0, C_s3_9_0;
FA FA_s3_9_0(.A_i(S_s4_9_2), .B_i(S_s4_9_1), .c_in(S_s4_9_0), .S_o(S_s3_9_0), .c_out(C_s3_9_0));
logic S_s3_9_1, C_s3_9_1;
FA FA_s3_9_1(.A_i(C_s4_8_2), .B_i(C_s4_8_1), .c_in(C_s4_8_0), .S_o(S_s3_9_1), .c_out(C_s3_9_1));
logic S_s3_10_0, C_s3_10_0;
FA FA_s3_10_0(.A_i(S_s4_10_2), .B_i(S_s4_10_1), .c_in(S_s4_10_0), .S_o(S_s3_10_0), .c_out(C_s3_10_0));
logic S_s3_10_1, C_s3_10_1;
FA FA_s3_10_1(.A_i(C_s4_9_2), .B_i(C_s4_9_1), .c_in(C_s4_9_0), .S_o(S_s3_10_1), .c_out(C_s3_10_1));
logic S_s3_11_0, C_s3_11_0;
FA FA_s3_11_0(.A_i(S_s4_11_2), .B_i(S_s4_11_1), .c_in(S_s4_11_0), .S_o(S_s3_11_0), .c_out(C_s3_11_0));
logic S_s3_11_1, C_s3_11_1;
FA FA_s3_11_1(.A_i(C_s4_10_2), .B_i(C_s4_10_1), .c_in(C_s4_10_0), .S_o(S_s3_11_1), .c_out(C_s3_11_1));
logic S_s3_12_0, C_s3_12_0;
FA FA_s3_12_0(.A_i(S_s4_12_2), .B_i(S_s4_12_1), .c_in(S_s4_12_0), .S_o(S_s3_12_0), .c_out(C_s3_12_0));
logic S_s3_12_1, C_s3_12_1;
FA FA_s3_12_1(.A_i(C_s4_11_2), .B_i(C_s4_11_1), .c_in(C_s4_11_0), .S_o(S_s3_12_1), .c_out(C_s3_12_1));
logic S_s3_13_0, C_s3_13_0;
FA FA_s3_13_0(.A_i(S_s4_13_2), .B_i(S_s4_13_1), .c_in(S_s4_13_0), .S_o(S_s3_13_0), .c_out(C_s3_13_0));
logic S_s3_13_1, C_s3_13_1;
FA FA_s3_13_1(.A_i(C_s4_12_2), .B_i(C_s4_12_1), .c_in(C_s4_12_0), .S_o(S_s3_13_1), .c_out(C_s3_13_1));
logic S_s3_14_0, C_s3_14_0;
FA FA_s3_14_0(.A_i(S_s4_14_2), .B_i(S_s4_14_1), .c_in(S_s4_14_0), .S_o(S_s3_14_0), .c_out(C_s3_14_0));
logic S_s3_14_1, C_s3_14_1;
FA FA_s3_14_1(.A_i(C_s4_13_2), .B_i(C_s4_13_1), .c_in(C_s4_13_0), .S_o(S_s3_14_1), .c_out(C_s3_14_1));
logic S_s3_15_0, C_s3_15_0;
FA FA_s3_15_0(.A_i(S_s4_15_2), .B_i(S_s4_15_1), .c_in(S_s4_15_0), .S_o(S_s3_15_0), .c_out(C_s3_15_0));
logic S_s3_15_1, C_s3_15_1;
FA FA_s3_15_1(.A_i(C_s4_14_2), .B_i(C_s4_14_1), .c_in(C_s4_14_0), .S_o(S_s3_15_1), .c_out(C_s3_15_1));
logic S_s3_16_0, C_s3_16_0;
FA FA_s3_16_0(.A_i(S_s4_16_2), .B_i(S_s4_16_1), .c_in(S_s4_16_0), .S_o(S_s3_16_0), .c_out(C_s3_16_0));
logic S_s3_16_1, C_s3_16_1;
FA FA_s3_16_1(.A_i(C_s4_15_2), .B_i(C_s4_15_1), .c_in(C_s4_15_0), .S_o(S_s3_16_1), .c_out(C_s3_16_1));
logic S_s3_17_0, C_s3_17_0;
FA FA_s3_17_0(.A_i(S_s4_17_2), .B_i(S_s4_17_1), .c_in(S_s4_17_0), .S_o(S_s3_17_0), .c_out(C_s3_17_0));
logic S_s3_17_1, C_s3_17_1;
FA FA_s3_17_1(.A_i(C_s4_16_2), .B_i(C_s4_16_1), .c_in(C_s4_16_0), .S_o(S_s3_17_1), .c_out(C_s3_17_1));
logic S_s3_18_0, C_s3_18_0;
FA FA_s3_18_0(.A_i(S_s4_18_2), .B_i(S_s4_18_1), .c_in(S_s4_18_0), .S_o(S_s3_18_0), .c_out(C_s3_18_0));
logic S_s3_18_1, C_s3_18_1;
FA FA_s3_18_1(.A_i(C_s4_17_2), .B_i(C_s4_17_1), .c_in(C_s4_17_0), .S_o(S_s3_18_1), .c_out(C_s3_18_1));
logic S_s3_19_0, C_s3_19_0;
FA FA_s3_19_0(.A_i(S_s4_19_2), .B_i(S_s4_19_1), .c_in(S_s4_19_0), .S_o(S_s3_19_0), .c_out(C_s3_19_0));
logic S_s3_19_1, C_s3_19_1;
FA FA_s3_19_1(.A_i(C_s4_18_2), .B_i(C_s4_18_1), .c_in(C_s4_18_0), .S_o(S_s3_19_1), .c_out(C_s3_19_1));
logic S_s3_20_0, C_s3_20_0;
FA FA_s3_20_0(.A_i(S_s4_20_2), .B_i(S_s4_20_1), .c_in(S_s4_20_0), .S_o(S_s3_20_0), .c_out(C_s3_20_0));
logic S_s3_20_1, C_s3_20_1;
FA FA_s3_20_1(.A_i(C_s4_19_2), .B_i(C_s4_19_1), .c_in(C_s4_19_0), .S_o(S_s3_20_1), .c_out(C_s3_20_1));
logic S_s3_21_0, C_s3_21_0;
FA FA_s3_21_0(.A_i(S_s4_21_2), .B_i(S_s4_21_1), .c_in(S_s4_21_0), .S_o(S_s3_21_0), .c_out(C_s3_21_0));
logic S_s3_21_1, C_s3_21_1;
FA FA_s3_21_1(.A_i(C_s4_20_2), .B_i(C_s4_20_1), .c_in(C_s4_20_0), .S_o(S_s3_21_1), .c_out(C_s3_21_1));
logic S_s3_22_0, C_s3_22_0;
FA FA_s3_22_0(.A_i(S_s4_22_2), .B_i(S_s4_22_1), .c_in(S_s4_22_0), .S_o(S_s3_22_0), .c_out(C_s3_22_0));
logic S_s3_22_1, C_s3_22_1;
FA FA_s3_22_1(.A_i(C_s4_21_2), .B_i(C_s4_21_1), .c_in(C_s4_21_0), .S_o(S_s3_22_1), .c_out(C_s3_22_1));
logic S_s3_23_0, C_s3_23_0;
FA FA_s3_23_0(.A_i(S_s4_23_2), .B_i(S_s4_23_1), .c_in(S_s4_23_0), .S_o(S_s3_23_0), .c_out(C_s3_23_0));
logic S_s3_23_1, C_s3_23_1;
FA FA_s3_23_1(.A_i(C_s4_22_2), .B_i(C_s4_22_1), .c_in(C_s4_22_0), .S_o(S_s3_23_1), .c_out(C_s3_23_1));
logic S_s3_24_0, C_s3_24_0;
FA FA_s3_24_0(.A_i(S_s4_24_2), .B_i(S_s4_24_1), .c_in(S_s4_24_0), .S_o(S_s3_24_0), .c_out(C_s3_24_0));
logic S_s3_24_1, C_s3_24_1;
FA FA_s3_24_1(.A_i(C_s4_23_2), .B_i(C_s4_23_1), .c_in(C_s4_23_0), .S_o(S_s3_24_1), .c_out(C_s3_24_1));
logic S_s3_25_0, C_s3_25_0;
FA FA_s3_25_0(.A_i(S_s4_25_2), .B_i(S_s4_25_1), .c_in(S_s4_25_0), .S_o(S_s3_25_0), .c_out(C_s3_25_0));
logic S_s3_25_1, C_s3_25_1;
FA FA_s3_25_1(.A_i(C_s4_24_2), .B_i(C_s4_24_1), .c_in(C_s4_24_0), .S_o(S_s3_25_1), .c_out(C_s3_25_1));
logic S_s3_26_0, C_s3_26_0;
FA FA_s3_26_0(.A_i(S_s4_26_2), .B_i(S_s4_26_1), .c_in(S_s4_26_0), .S_o(S_s3_26_0), .c_out(C_s3_26_0));
logic S_s3_26_1, C_s3_26_1;
FA FA_s3_26_1(.A_i(C_s4_25_2), .B_i(C_s4_25_1), .c_in(C_s4_25_0), .S_o(S_s3_26_1), .c_out(C_s3_26_1));
logic S_s3_27_0, C_s3_27_0;
FA FA_s3_27_0(.A_i(S_s4_27_2), .B_i(S_s4_27_1), .c_in(S_s4_27_0), .S_o(S_s3_27_0), .c_out(C_s3_27_0));
logic S_s3_27_1, C_s3_27_1;
FA FA_s3_27_1(.A_i(C_s4_26_2), .B_i(C_s4_26_1), .c_in(C_s4_26_0), .S_o(S_s3_27_1), .c_out(C_s3_27_1));
logic S_s3_28_0, C_s3_28_0;
FA FA_s3_28_0(.A_i(S_s4_28_2), .B_i(S_s4_28_1), .c_in(S_s4_28_0), .S_o(S_s3_28_0), .c_out(C_s3_28_0));
logic S_s3_28_1, C_s3_28_1;
FA FA_s3_28_1(.A_i(C_s4_27_2), .B_i(C_s4_27_1), .c_in(C_s4_27_0), .S_o(S_s3_28_1), .c_out(C_s3_28_1));
logic S_s3_29_0, C_s3_29_0;
FA FA_s3_29_0(.A_i(S_s4_29_2), .B_i(S_s4_29_1), .c_in(S_s4_29_0), .S_o(S_s3_29_0), .c_out(C_s3_29_0));
logic S_s3_29_1, C_s3_29_1;
FA FA_s3_29_1(.A_i(C_s4_28_2), .B_i(C_s4_28_1), .c_in(C_s4_28_0), .S_o(S_s3_29_1), .c_out(C_s3_29_1));
logic S_s3_30_0, C_s3_30_0;
FA FA_s3_30_0(.A_i(S_s4_30_2), .B_i(S_s4_30_1), .c_in(S_s4_30_0), .S_o(S_s3_30_0), .c_out(C_s3_30_0));
logic S_s3_30_1, C_s3_30_1;
FA FA_s3_30_1(.A_i(C_s4_29_2), .B_i(C_s4_29_1), .c_in(C_s4_29_0), .S_o(S_s3_30_1), .c_out(C_s3_30_1));
logic S_s3_31_0, C_s3_31_0;
FA FA_s3_31_0(.A_i(S_s4_31_2), .B_i(S_s4_31_1), .c_in(S_s4_31_0), .S_o(S_s3_31_0), .c_out(C_s3_31_0));
logic S_s3_31_1, C_s3_31_1;
FA FA_s3_31_1(.A_i(C_s4_30_2), .B_i(C_s4_30_1), .c_in(C_s4_30_0), .S_o(S_s3_31_1), .c_out(C_s3_31_1));
logic S_s3_32_0, C_s3_32_0;
FA FA_s3_32_0(.A_i(S_s4_32_2), .B_i(S_s4_32_1), .c_in(S_s4_32_0), .S_o(S_s3_32_0), .c_out(C_s3_32_0));
logic S_s3_32_1, C_s3_32_1;
FA FA_s3_32_1(.A_i(C_s4_31_2), .B_i(C_s4_31_1), .c_in(C_s4_31_0), .S_o(S_s3_32_1), .c_out(C_s3_32_1));
logic S_s3_33_0, C_s3_33_0;
FA FA_s3_33_0(.A_i(S_s4_33_2), .B_i(S_s4_33_1), .c_in(S_s4_33_0), .S_o(S_s3_33_0), .c_out(C_s3_33_0));
logic S_s3_33_1, C_s3_33_1;
FA FA_s3_33_1(.A_i(C_s4_32_2), .B_i(C_s4_32_1), .c_in(C_s4_32_0), .S_o(S_s3_33_1), .c_out(C_s3_33_1));
logic S_s3_34_0, C_s3_34_0;
FA FA_s3_34_0(.A_i(S_s4_34_2), .B_i(S_s4_34_1), .c_in(S_s4_34_0), .S_o(S_s3_34_0), .c_out(C_s3_34_0));
logic S_s3_34_1, C_s3_34_1;
FA FA_s3_34_1(.A_i(C_s4_33_2), .B_i(C_s4_33_1), .c_in(C_s4_33_0), .S_o(S_s3_34_1), .c_out(C_s3_34_1));
logic S_s3_35_0, C_s3_35_0;
FA FA_s3_35_0(.A_i(S_s4_35_2), .B_i(S_s4_35_1), .c_in(S_s4_35_0), .S_o(S_s3_35_0), .c_out(C_s3_35_0));
logic S_s3_35_1, C_s3_35_1;
FA FA_s3_35_1(.A_i(C_s4_34_2), .B_i(C_s4_34_1), .c_in(C_s4_34_0), .S_o(S_s3_35_1), .c_out(C_s3_35_1));
logic S_s3_36_0, C_s3_36_0;
FA FA_s3_36_0(.A_i(S_s4_36_2), .B_i(S_s4_36_1), .c_in(S_s4_36_0), .S_o(S_s3_36_0), .c_out(C_s3_36_0));
logic S_s3_36_1, C_s3_36_1;
FA FA_s3_36_1(.A_i(C_s4_35_2), .B_i(C_s4_35_1), .c_in(C_s4_35_0), .S_o(S_s3_36_1), .c_out(C_s3_36_1));
logic S_s3_37_0, C_s3_37_0;
FA FA_s3_37_0(.A_i(S_s4_37_2), .B_i(S_s4_37_1), .c_in(S_s4_37_0), .S_o(S_s3_37_0), .c_out(C_s3_37_0));
logic S_s3_37_1, C_s3_37_1;
FA FA_s3_37_1(.A_i(C_s4_36_2), .B_i(C_s4_36_1), .c_in(C_s4_36_0), .S_o(S_s3_37_1), .c_out(C_s3_37_1));
logic S_s3_38_0, C_s3_38_0;
FA FA_s3_38_0(.A_i(S_s4_38_2), .B_i(S_s4_38_1), .c_in(S_s4_38_0), .S_o(S_s3_38_0), .c_out(C_s3_38_0));
logic S_s3_38_1, C_s3_38_1;
FA FA_s3_38_1(.A_i(C_s4_37_2), .B_i(C_s4_37_1), .c_in(C_s4_37_0), .S_o(S_s3_38_1), .c_out(C_s3_38_1));
logic S_s3_39_0, C_s3_39_0;
FA FA_s3_39_0(.A_i(S_s4_39_2), .B_i(S_s4_39_1), .c_in(S_s4_39_0), .S_o(S_s3_39_0), .c_out(C_s3_39_0));
logic S_s3_39_1, C_s3_39_1;
FA FA_s3_39_1(.A_i(C_s4_38_2), .B_i(C_s4_38_1), .c_in(C_s4_38_0), .S_o(S_s3_39_1), .c_out(C_s3_39_1));
logic S_s3_40_0, C_s3_40_0;
FA FA_s3_40_0(.A_i(S_s4_40_2), .B_i(S_s4_40_1), .c_in(S_s4_40_0), .S_o(S_s3_40_0), .c_out(C_s3_40_0));
logic S_s3_40_1, C_s3_40_1;
FA FA_s3_40_1(.A_i(C_s4_39_2), .B_i(C_s4_39_1), .c_in(C_s4_39_0), .S_o(S_s3_40_1), .c_out(C_s3_40_1));
logic S_s3_41_0, C_s3_41_0;
FA FA_s3_41_0(.A_i(S_s4_41_2), .B_i(S_s4_41_1), .c_in(S_s4_41_0), .S_o(S_s3_41_0), .c_out(C_s3_41_0));
logic S_s3_41_1, C_s3_41_1;
FA FA_s3_41_1(.A_i(C_s4_40_2), .B_i(C_s4_40_1), .c_in(C_s4_40_0), .S_o(S_s3_41_1), .c_out(C_s3_41_1));
logic S_s3_42_0, C_s3_42_0;
FA FA_s3_42_0(.A_i(S_s4_42_2), .B_i(S_s4_42_1), .c_in(S_s4_42_0), .S_o(S_s3_42_0), .c_out(C_s3_42_0));
logic S_s3_42_1, C_s3_42_1;
FA FA_s3_42_1(.A_i(C_s4_41_2), .B_i(C_s4_41_1), .c_in(C_s4_41_0), .S_o(S_s3_42_1), .c_out(C_s3_42_1));
logic S_s3_43_0, C_s3_43_0;
FA FA_s3_43_0(.A_i(S_s4_43_2), .B_i(S_s4_43_1), .c_in(S_s4_43_0), .S_o(S_s3_43_0), .c_out(C_s3_43_0));
logic S_s3_43_1, C_s3_43_1;
FA FA_s3_43_1(.A_i(C_s4_42_2), .B_i(C_s4_42_1), .c_in(C_s4_42_0), .S_o(S_s3_43_1), .c_out(C_s3_43_1));
logic S_s3_44_0, C_s3_44_0;
FA FA_s3_44_0(.A_i(S_s4_44_2), .B_i(S_s4_44_1), .c_in(S_s4_44_0), .S_o(S_s3_44_0), .c_out(C_s3_44_0));
logic S_s3_44_1, C_s3_44_1;
FA FA_s3_44_1(.A_i(C_s4_43_2), .B_i(C_s4_43_1), .c_in(C_s4_43_0), .S_o(S_s3_44_1), .c_out(C_s3_44_1));
logic S_s3_45_0, C_s3_45_0;
FA FA_s3_45_0(.A_i(S_s4_45_2), .B_i(S_s4_45_1), .c_in(S_s4_45_0), .S_o(S_s3_45_0), .c_out(C_s3_45_0));
logic S_s3_45_1, C_s3_45_1;
FA FA_s3_45_1(.A_i(C_s4_44_2), .B_i(C_s4_44_1), .c_in(C_s4_44_0), .S_o(S_s3_45_1), .c_out(C_s3_45_1));
logic S_s3_46_0, C_s3_46_0;
FA FA_s3_46_0(.A_i(S_s4_46_2), .B_i(S_s4_46_1), .c_in(S_s4_46_0), .S_o(S_s3_46_0), .c_out(C_s3_46_0));
logic S_s3_46_1, C_s3_46_1;
FA FA_s3_46_1(.A_i(C_s4_45_2), .B_i(C_s4_45_1), .c_in(C_s4_45_0), .S_o(S_s3_46_1), .c_out(C_s3_46_1));
logic S_s3_47_0, C_s3_47_0;
FA FA_s3_47_0(.A_i(S_s4_47_2), .B_i(S_s4_47_1), .c_in(S_s4_47_0), .S_o(S_s3_47_0), .c_out(C_s3_47_0));
logic S_s3_47_1, C_s3_47_1;
FA FA_s3_47_1(.A_i(C_s4_46_2), .B_i(C_s4_46_1), .c_in(C_s4_46_0), .S_o(S_s3_47_1), .c_out(C_s3_47_1));
logic S_s3_48_0, C_s3_48_0;
FA FA_s3_48_0(.A_i(S_s4_48_2), .B_i(S_s4_48_1), .c_in(S_s4_48_0), .S_o(S_s3_48_0), .c_out(C_s3_48_0));
logic S_s3_48_1, C_s3_48_1;
FA FA_s3_48_1(.A_i(C_s4_47_2), .B_i(C_s4_47_1), .c_in(C_s4_47_0), .S_o(S_s3_48_1), .c_out(C_s3_48_1));
logic S_s3_49_0, C_s3_49_0;
FA FA_s3_49_0(.A_i(S_s4_49_2), .B_i(S_s4_49_1), .c_in(S_s4_49_0), .S_o(S_s3_49_0), .c_out(C_s3_49_0));
logic S_s3_49_1, C_s3_49_1;
FA FA_s3_49_1(.A_i(C_s4_48_2), .B_i(C_s4_48_1), .c_in(C_s4_48_0), .S_o(S_s3_49_1), .c_out(C_s3_49_1));
logic S_s3_50_0, C_s3_50_0;
FA FA_s3_50_0(.A_i(S_s4_50_2), .B_i(S_s4_50_1), .c_in(S_s4_50_0), .S_o(S_s3_50_0), .c_out(C_s3_50_0));
logic S_s3_50_1, C_s3_50_1;
FA FA_s3_50_1(.A_i(C_s4_49_2), .B_i(C_s4_49_1), .c_in(C_s4_49_0), .S_o(S_s3_50_1), .c_out(C_s3_50_1));
logic S_s3_51_0, C_s3_51_0;
FA FA_s3_51_0(.A_i(S_s4_51_2), .B_i(S_s4_51_1), .c_in(S_s4_51_0), .S_o(S_s3_51_0), .c_out(C_s3_51_0));
logic S_s3_51_1, C_s3_51_1;
FA FA_s3_51_1(.A_i(C_s4_50_2), .B_i(C_s4_50_1), .c_in(C_s4_50_0), .S_o(S_s3_51_1), .c_out(C_s3_51_1));
logic S_s3_52_0, C_s3_52_0;
FA FA_s3_52_0(.A_i(S_s4_52_2), .B_i(S_s4_52_1), .c_in(S_s4_52_0), .S_o(S_s3_52_0), .c_out(C_s3_52_0));
logic S_s3_52_1, C_s3_52_1;
FA FA_s3_52_1(.A_i(C_s4_51_2), .B_i(C_s4_51_1), .c_in(C_s4_51_0), .S_o(S_s3_52_1), .c_out(C_s3_52_1));
logic S_s3_53_0, C_s3_53_0;
FA FA_s3_53_0(.A_i(S_s4_53_2), .B_i(S_s4_53_1), .c_in(S_s4_53_0), .S_o(S_s3_53_0), .c_out(C_s3_53_0));
logic S_s3_53_1, C_s3_53_1;
FA FA_s3_53_1(.A_i(C_s4_52_2), .B_i(C_s4_52_1), .c_in(C_s4_52_0), .S_o(S_s3_53_1), .c_out(C_s3_53_1));
logic S_s3_54_0, C_s3_54_0;
FA FA_s3_54_0(.A_i(S_s4_54_2), .B_i(S_s4_54_1), .c_in(S_s4_54_0), .S_o(S_s3_54_0), .c_out(C_s3_54_0));
logic S_s3_54_1, C_s3_54_1;
FA FA_s3_54_1(.A_i(C_s4_53_2), .B_i(C_s4_53_1), .c_in(C_s4_53_0), .S_o(S_s3_54_1), .c_out(C_s3_54_1));
logic S_s3_55_0, C_s3_55_0;
FA FA_s3_55_0(.A_i(S_s4_55_2), .B_i(S_s4_55_1), .c_in(S_s4_55_0), .S_o(S_s3_55_0), .c_out(C_s3_55_0));
logic S_s3_55_1, C_s3_55_1;
FA FA_s3_55_1(.A_i(C_s4_54_2), .B_i(C_s4_54_1), .c_in(C_s4_54_0), .S_o(S_s3_55_1), .c_out(C_s3_55_1));
logic S_s3_56_0, C_s3_56_0;
FA FA_s3_56_0(.A_i(S_s4_56_1), .B_i(S_s4_56_0), .c_in(C_s4_55_2), .S_o(S_s3_56_0), .c_out(C_s3_56_0));
logic S_s3_56_1, C_s3_56_1;
FA FA_s3_56_1(.A_i(C_s4_55_1), .B_i(C_s4_55_0), .c_in(comb[31][25]), .S_o(S_s3_56_1), .c_out(C_s3_56_1));
logic S_s3_57_0, C_s3_57_0;
FA FA_s3_57_0(.A_i(S_s4_57_0), .B_i(C_s4_56_1), .c_in(C_s4_56_0), .S_o(S_s3_57_0), .c_out(C_s3_57_0));
logic S_s3_57_1, C_s3_57_1;
FA FA_s3_57_1(.A_i(comb[29][28]), .B_i(comb[30][27]), .c_in(comb[31][26]), .S_o(S_s3_57_1), .c_out(C_s3_57_1));
logic S_s3_58_0, C_s3_58_0;
FA FA_s3_58_0(.A_i(C_s4_57_0), .B_i(comb[27][31]), .c_in(comb[28][30]), .S_o(S_s3_58_0), .c_out(C_s3_58_0));
logic S_s3_58_1, C_s3_58_1;
FA FA_s3_58_1(.A_i(comb[29][29]), .B_i(comb[30][28]), .c_in(comb[31][27]), .S_o(S_s3_58_1), .c_out(C_s3_58_1));
logic S_s3_59_0, C_s3_59_0;
FA FA_s3_59_0(.A_i(comb[28][31]), .B_i(comb[29][30]), .c_in(comb[30][29]), .S_o(S_s3_59_0), .c_out(C_s3_59_0));
// stage 3 end ======================================================================================================= 

// stage 2 begin ======================================================================================================= 
logic S_s2_3_0, C_s2_3_0;
HA HA_s2_30(.A_i(comb[0][3]), .B_i(comb[1][2]), .S_o(S_s2_3_0), .c_out(C_s2_3_0));
logic S_s2_4_0, C_s2_4_0;
FA FA_s2_4_0(.A_i(S_s3_4_0), .B_i(comb[2][2]), .c_in(comb[3][1]), .S_o(S_s2_4_0), .c_out(C_s2_4_0));
logic S_s2_5_0, C_s2_5_0;
FA FA_s2_5_0(.A_i(S_s3_5_1), .B_i(S_s3_5_0), .c_in(C_s3_4_0), .S_o(S_s2_5_0), .c_out(C_s2_5_0));
logic S_s2_6_0, C_s2_6_0;
FA FA_s2_6_0(.A_i(S_s3_6_1), .B_i(S_s3_6_0), .c_in(C_s3_5_1), .S_o(S_s2_6_0), .c_out(C_s2_6_0));
logic S_s2_7_0, C_s2_7_0;
FA FA_s2_7_0(.A_i(S_s3_7_1), .B_i(S_s3_7_0), .c_in(C_s3_6_1), .S_o(S_s2_7_0), .c_out(C_s2_7_0));
logic S_s2_8_0, C_s2_8_0;
FA FA_s2_8_0(.A_i(S_s3_8_1), .B_i(S_s3_8_0), .c_in(C_s3_7_1), .S_o(S_s2_8_0), .c_out(C_s2_8_0));
logic S_s2_9_0, C_s2_9_0;
FA FA_s2_9_0(.A_i(S_s3_9_1), .B_i(S_s3_9_0), .c_in(C_s3_8_1), .S_o(S_s2_9_0), .c_out(C_s2_9_0));
logic S_s2_10_0, C_s2_10_0;
FA FA_s2_10_0(.A_i(S_s3_10_1), .B_i(S_s3_10_0), .c_in(C_s3_9_1), .S_o(S_s2_10_0), .c_out(C_s2_10_0));
logic S_s2_11_0, C_s2_11_0;
FA FA_s2_11_0(.A_i(S_s3_11_1), .B_i(S_s3_11_0), .c_in(C_s3_10_1), .S_o(S_s2_11_0), .c_out(C_s2_11_0));
logic S_s2_12_0, C_s2_12_0;
FA FA_s2_12_0(.A_i(S_s3_12_1), .B_i(S_s3_12_0), .c_in(C_s3_11_1), .S_o(S_s2_12_0), .c_out(C_s2_12_0));
logic S_s2_13_0, C_s2_13_0;
FA FA_s2_13_0(.A_i(S_s3_13_1), .B_i(S_s3_13_0), .c_in(C_s3_12_1), .S_o(S_s2_13_0), .c_out(C_s2_13_0));
logic S_s2_14_0, C_s2_14_0;
FA FA_s2_14_0(.A_i(S_s3_14_1), .B_i(S_s3_14_0), .c_in(C_s3_13_1), .S_o(S_s2_14_0), .c_out(C_s2_14_0));
logic S_s2_15_0, C_s2_15_0;
FA FA_s2_15_0(.A_i(S_s3_15_1), .B_i(S_s3_15_0), .c_in(C_s3_14_1), .S_o(S_s2_15_0), .c_out(C_s2_15_0));
logic S_s2_16_0, C_s2_16_0;
FA FA_s2_16_0(.A_i(S_s3_16_1), .B_i(S_s3_16_0), .c_in(C_s3_15_1), .S_o(S_s2_16_0), .c_out(C_s2_16_0));
logic S_s2_17_0, C_s2_17_0;
FA FA_s2_17_0(.A_i(S_s3_17_1), .B_i(S_s3_17_0), .c_in(C_s3_16_1), .S_o(S_s2_17_0), .c_out(C_s2_17_0));
logic S_s2_18_0, C_s2_18_0;
FA FA_s2_18_0(.A_i(S_s3_18_1), .B_i(S_s3_18_0), .c_in(C_s3_17_1), .S_o(S_s2_18_0), .c_out(C_s2_18_0));
logic S_s2_19_0, C_s2_19_0;
FA FA_s2_19_0(.A_i(S_s3_19_1), .B_i(S_s3_19_0), .c_in(C_s3_18_1), .S_o(S_s2_19_0), .c_out(C_s2_19_0));
logic S_s2_20_0, C_s2_20_0;
FA FA_s2_20_0(.A_i(S_s3_20_1), .B_i(S_s3_20_0), .c_in(C_s3_19_1), .S_o(S_s2_20_0), .c_out(C_s2_20_0));
logic S_s2_21_0, C_s2_21_0;
FA FA_s2_21_0(.A_i(S_s3_21_1), .B_i(S_s3_21_0), .c_in(C_s3_20_1), .S_o(S_s2_21_0), .c_out(C_s2_21_0));
logic S_s2_22_0, C_s2_22_0;
FA FA_s2_22_0(.A_i(S_s3_22_1), .B_i(S_s3_22_0), .c_in(C_s3_21_1), .S_o(S_s2_22_0), .c_out(C_s2_22_0));
logic S_s2_23_0, C_s2_23_0;
FA FA_s2_23_0(.A_i(S_s3_23_1), .B_i(S_s3_23_0), .c_in(C_s3_22_1), .S_o(S_s2_23_0), .c_out(C_s2_23_0));
logic S_s2_24_0, C_s2_24_0;
FA FA_s2_24_0(.A_i(S_s3_24_1), .B_i(S_s3_24_0), .c_in(C_s3_23_1), .S_o(S_s2_24_0), .c_out(C_s2_24_0));
logic S_s2_25_0, C_s2_25_0;
FA FA_s2_25_0(.A_i(S_s3_25_1), .B_i(S_s3_25_0), .c_in(C_s3_24_1), .S_o(S_s2_25_0), .c_out(C_s2_25_0));
logic S_s2_26_0, C_s2_26_0;
FA FA_s2_26_0(.A_i(S_s3_26_1), .B_i(S_s3_26_0), .c_in(C_s3_25_1), .S_o(S_s2_26_0), .c_out(C_s2_26_0));
logic S_s2_27_0, C_s2_27_0;
FA FA_s2_27_0(.A_i(S_s3_27_1), .B_i(S_s3_27_0), .c_in(C_s3_26_1), .S_o(S_s2_27_0), .c_out(C_s2_27_0));
logic S_s2_28_0, C_s2_28_0;
FA FA_s2_28_0(.A_i(S_s3_28_1), .B_i(S_s3_28_0), .c_in(C_s3_27_1), .S_o(S_s2_28_0), .c_out(C_s2_28_0));
logic S_s2_29_0, C_s2_29_0;
FA FA_s2_29_0(.A_i(S_s3_29_1), .B_i(S_s3_29_0), .c_in(C_s3_28_1), .S_o(S_s2_29_0), .c_out(C_s2_29_0));
logic S_s2_30_0, C_s2_30_0;
FA FA_s2_30_0(.A_i(S_s3_30_1), .B_i(S_s3_30_0), .c_in(C_s3_29_1), .S_o(S_s2_30_0), .c_out(C_s2_30_0));
logic S_s2_31_0, C_s2_31_0;
FA FA_s2_31_0(.A_i(S_s3_31_1), .B_i(S_s3_31_0), .c_in(C_s3_30_1), .S_o(S_s2_31_0), .c_out(C_s2_31_0));
logic S_s2_32_0, C_s2_32_0;
FA FA_s2_32_0(.A_i(S_s3_32_1), .B_i(S_s3_32_0), .c_in(C_s3_31_1), .S_o(S_s2_32_0), .c_out(C_s2_32_0));
logic S_s2_33_0, C_s2_33_0;
FA FA_s2_33_0(.A_i(S_s3_33_1), .B_i(S_s3_33_0), .c_in(C_s3_32_1), .S_o(S_s2_33_0), .c_out(C_s2_33_0));
logic S_s2_34_0, C_s2_34_0;
FA FA_s2_34_0(.A_i(S_s3_34_1), .B_i(S_s3_34_0), .c_in(C_s3_33_1), .S_o(S_s2_34_0), .c_out(C_s2_34_0));
logic S_s2_35_0, C_s2_35_0;
FA FA_s2_35_0(.A_i(S_s3_35_1), .B_i(S_s3_35_0), .c_in(C_s3_34_1), .S_o(S_s2_35_0), .c_out(C_s2_35_0));
logic S_s2_36_0, C_s2_36_0;
FA FA_s2_36_0(.A_i(S_s3_36_1), .B_i(S_s3_36_0), .c_in(C_s3_35_1), .S_o(S_s2_36_0), .c_out(C_s2_36_0));
logic S_s2_37_0, C_s2_37_0;
FA FA_s2_37_0(.A_i(S_s3_37_1), .B_i(S_s3_37_0), .c_in(C_s3_36_1), .S_o(S_s2_37_0), .c_out(C_s2_37_0));
logic S_s2_38_0, C_s2_38_0;
FA FA_s2_38_0(.A_i(S_s3_38_1), .B_i(S_s3_38_0), .c_in(C_s3_37_1), .S_o(S_s2_38_0), .c_out(C_s2_38_0));
logic S_s2_39_0, C_s2_39_0;
FA FA_s2_39_0(.A_i(S_s3_39_1), .B_i(S_s3_39_0), .c_in(C_s3_38_1), .S_o(S_s2_39_0), .c_out(C_s2_39_0));
logic S_s2_40_0, C_s2_40_0;
FA FA_s2_40_0(.A_i(S_s3_40_1), .B_i(S_s3_40_0), .c_in(C_s3_39_1), .S_o(S_s2_40_0), .c_out(C_s2_40_0));
logic S_s2_41_0, C_s2_41_0;
FA FA_s2_41_0(.A_i(S_s3_41_1), .B_i(S_s3_41_0), .c_in(C_s3_40_1), .S_o(S_s2_41_0), .c_out(C_s2_41_0));
logic S_s2_42_0, C_s2_42_0;
FA FA_s2_42_0(.A_i(S_s3_42_1), .B_i(S_s3_42_0), .c_in(C_s3_41_1), .S_o(S_s2_42_0), .c_out(C_s2_42_0));
logic S_s2_43_0, C_s2_43_0;
FA FA_s2_43_0(.A_i(S_s3_43_1), .B_i(S_s3_43_0), .c_in(C_s3_42_1), .S_o(S_s2_43_0), .c_out(C_s2_43_0));
logic S_s2_44_0, C_s2_44_0;
FA FA_s2_44_0(.A_i(S_s3_44_1), .B_i(S_s3_44_0), .c_in(C_s3_43_1), .S_o(S_s2_44_0), .c_out(C_s2_44_0));
logic S_s2_45_0, C_s2_45_0;
FA FA_s2_45_0(.A_i(S_s3_45_1), .B_i(S_s3_45_0), .c_in(C_s3_44_1), .S_o(S_s2_45_0), .c_out(C_s2_45_0));
logic S_s2_46_0, C_s2_46_0;
FA FA_s2_46_0(.A_i(S_s3_46_1), .B_i(S_s3_46_0), .c_in(C_s3_45_1), .S_o(S_s2_46_0), .c_out(C_s2_46_0));
logic S_s2_47_0, C_s2_47_0;
FA FA_s2_47_0(.A_i(S_s3_47_1), .B_i(S_s3_47_0), .c_in(C_s3_46_1), .S_o(S_s2_47_0), .c_out(C_s2_47_0));
logic S_s2_48_0, C_s2_48_0;
FA FA_s2_48_0(.A_i(S_s3_48_1), .B_i(S_s3_48_0), .c_in(C_s3_47_1), .S_o(S_s2_48_0), .c_out(C_s2_48_0));
logic S_s2_49_0, C_s2_49_0;
FA FA_s2_49_0(.A_i(S_s3_49_1), .B_i(S_s3_49_0), .c_in(C_s3_48_1), .S_o(S_s2_49_0), .c_out(C_s2_49_0));
logic S_s2_50_0, C_s2_50_0;
FA FA_s2_50_0(.A_i(S_s3_50_1), .B_i(S_s3_50_0), .c_in(C_s3_49_1), .S_o(S_s2_50_0), .c_out(C_s2_50_0));
logic S_s2_51_0, C_s2_51_0;
FA FA_s2_51_0(.A_i(S_s3_51_1), .B_i(S_s3_51_0), .c_in(C_s3_50_1), .S_o(S_s2_51_0), .c_out(C_s2_51_0));
logic S_s2_52_0, C_s2_52_0;
FA FA_s2_52_0(.A_i(S_s3_52_1), .B_i(S_s3_52_0), .c_in(C_s3_51_1), .S_o(S_s2_52_0), .c_out(C_s2_52_0));
logic S_s2_53_0, C_s2_53_0;
FA FA_s2_53_0(.A_i(S_s3_53_1), .B_i(S_s3_53_0), .c_in(C_s3_52_1), .S_o(S_s2_53_0), .c_out(C_s2_53_0));
logic S_s2_54_0, C_s2_54_0;
FA FA_s2_54_0(.A_i(S_s3_54_1), .B_i(S_s3_54_0), .c_in(C_s3_53_1), .S_o(S_s2_54_0), .c_out(C_s2_54_0));
logic S_s2_55_0, C_s2_55_0;
FA FA_s2_55_0(.A_i(S_s3_55_1), .B_i(S_s3_55_0), .c_in(C_s3_54_1), .S_o(S_s2_55_0), .c_out(C_s2_55_0));
logic S_s2_56_0, C_s2_56_0;
FA FA_s2_56_0(.A_i(S_s3_56_1), .B_i(S_s3_56_0), .c_in(C_s3_55_1), .S_o(S_s2_56_0), .c_out(C_s2_56_0));
logic S_s2_57_0, C_s2_57_0;
FA FA_s2_57_0(.A_i(S_s3_57_1), .B_i(S_s3_57_0), .c_in(C_s3_56_1), .S_o(S_s2_57_0), .c_out(C_s2_57_0));
logic S_s2_58_0, C_s2_58_0;
FA FA_s2_58_0(.A_i(S_s3_58_1), .B_i(S_s3_58_0), .c_in(C_s3_57_1), .S_o(S_s2_58_0), .c_out(C_s2_58_0));
logic S_s2_59_0, C_s2_59_0;
FA FA_s2_59_0(.A_i(S_s3_59_0), .B_i(C_s3_58_1), .c_in(C_s3_58_0), .S_o(S_s2_59_0), .c_out(C_s2_59_0));
logic S_s2_60_0, C_s2_60_0;
FA FA_s2_60_0(.A_i(C_s3_59_0), .B_i(comb[29][31]), .c_in(comb[30][30]), .S_o(S_s2_60_0), .c_out(C_s2_60_0));
// stage 2 end ======================================================================================================= 

// stage 1 begin ======================================================================================================= 
logic S_s1_2_0, C_s1_2_0;
HA HA_s1_20(.A_i(comb[0][2]), .B_i(comb[1][1]), .S_o(S_s1_2_0), .c_out(C_s1_2_0));
logic S_s1_3_0, C_s1_3_0;
FA FA_s1_3_0(.A_i(S_s2_3_0), .B_i(comb[2][1]), .c_in(comb[3][0]), .S_o(S_s1_3_0), .c_out(C_s1_3_0));
logic S_s1_4_0, C_s1_4_0;
FA FA_s1_4_0(.A_i(S_s2_4_0), .B_i(C_s2_3_0), .c_in(comb[4][0]), .S_o(S_s1_4_0), .c_out(C_s1_4_0));
logic S_s1_5_0, C_s1_5_0;
FA FA_s1_5_0(.A_i(S_s2_5_0), .B_i(C_s2_4_0), .c_in(comb[5][0]), .S_o(S_s1_5_0), .c_out(C_s1_5_0));
logic S_s1_6_0, C_s1_6_0;
FA FA_s1_6_0(.A_i(S_s2_6_0), .B_i(C_s2_5_0), .c_in(C_s3_5_0), .S_o(S_s1_6_0), .c_out(C_s1_6_0));
logic S_s1_7_0, C_s1_7_0;
FA FA_s1_7_0(.A_i(S_s2_7_0), .B_i(C_s2_6_0), .c_in(C_s3_6_0), .S_o(S_s1_7_0), .c_out(C_s1_7_0));
logic S_s1_8_0, C_s1_8_0;
FA FA_s1_8_0(.A_i(S_s2_8_0), .B_i(C_s2_7_0), .c_in(C_s3_7_0), .S_o(S_s1_8_0), .c_out(C_s1_8_0));
logic S_s1_9_0, C_s1_9_0;
FA FA_s1_9_0(.A_i(S_s2_9_0), .B_i(C_s2_8_0), .c_in(C_s3_8_0), .S_o(S_s1_9_0), .c_out(C_s1_9_0));
logic S_s1_10_0, C_s1_10_0;
FA FA_s1_10_0(.A_i(S_s2_10_0), .B_i(C_s2_9_0), .c_in(C_s3_9_0), .S_o(S_s1_10_0), .c_out(C_s1_10_0));
logic S_s1_11_0, C_s1_11_0;
FA FA_s1_11_0(.A_i(S_s2_11_0), .B_i(C_s2_10_0), .c_in(C_s3_10_0), .S_o(S_s1_11_0), .c_out(C_s1_11_0));
logic S_s1_12_0, C_s1_12_0;
FA FA_s1_12_0(.A_i(S_s2_12_0), .B_i(C_s2_11_0), .c_in(C_s3_11_0), .S_o(S_s1_12_0), .c_out(C_s1_12_0));
logic S_s1_13_0, C_s1_13_0;
FA FA_s1_13_0(.A_i(S_s2_13_0), .B_i(C_s2_12_0), .c_in(C_s3_12_0), .S_o(S_s1_13_0), .c_out(C_s1_13_0));
logic S_s1_14_0, C_s1_14_0;
FA FA_s1_14_0(.A_i(S_s2_14_0), .B_i(C_s2_13_0), .c_in(C_s3_13_0), .S_o(S_s1_14_0), .c_out(C_s1_14_0));
logic S_s1_15_0, C_s1_15_0;
FA FA_s1_15_0(.A_i(S_s2_15_0), .B_i(C_s2_14_0), .c_in(C_s3_14_0), .S_o(S_s1_15_0), .c_out(C_s1_15_0));
logic S_s1_16_0, C_s1_16_0;
FA FA_s1_16_0(.A_i(S_s2_16_0), .B_i(C_s2_15_0), .c_in(C_s3_15_0), .S_o(S_s1_16_0), .c_out(C_s1_16_0));
logic S_s1_17_0, C_s1_17_0;
FA FA_s1_17_0(.A_i(S_s2_17_0), .B_i(C_s2_16_0), .c_in(C_s3_16_0), .S_o(S_s1_17_0), .c_out(C_s1_17_0));
logic S_s1_18_0, C_s1_18_0;
FA FA_s1_18_0(.A_i(S_s2_18_0), .B_i(C_s2_17_0), .c_in(C_s3_17_0), .S_o(S_s1_18_0), .c_out(C_s1_18_0));
logic S_s1_19_0, C_s1_19_0;
FA FA_s1_19_0(.A_i(S_s2_19_0), .B_i(C_s2_18_0), .c_in(C_s3_18_0), .S_o(S_s1_19_0), .c_out(C_s1_19_0));
logic S_s1_20_0, C_s1_20_0;
FA FA_s1_20_0(.A_i(S_s2_20_0), .B_i(C_s2_19_0), .c_in(C_s3_19_0), .S_o(S_s1_20_0), .c_out(C_s1_20_0));
logic S_s1_21_0, C_s1_21_0;
FA FA_s1_21_0(.A_i(S_s2_21_0), .B_i(C_s2_20_0), .c_in(C_s3_20_0), .S_o(S_s1_21_0), .c_out(C_s1_21_0));
logic S_s1_22_0, C_s1_22_0;
FA FA_s1_22_0(.A_i(S_s2_22_0), .B_i(C_s2_21_0), .c_in(C_s3_21_0), .S_o(S_s1_22_0), .c_out(C_s1_22_0));
logic S_s1_23_0, C_s1_23_0;
FA FA_s1_23_0(.A_i(S_s2_23_0), .B_i(C_s2_22_0), .c_in(C_s3_22_0), .S_o(S_s1_23_0), .c_out(C_s1_23_0));
logic S_s1_24_0, C_s1_24_0;
FA FA_s1_24_0(.A_i(S_s2_24_0), .B_i(C_s2_23_0), .c_in(C_s3_23_0), .S_o(S_s1_24_0), .c_out(C_s1_24_0));
logic S_s1_25_0, C_s1_25_0;
FA FA_s1_25_0(.A_i(S_s2_25_0), .B_i(C_s2_24_0), .c_in(C_s3_24_0), .S_o(S_s1_25_0), .c_out(C_s1_25_0));
logic S_s1_26_0, C_s1_26_0;
FA FA_s1_26_0(.A_i(S_s2_26_0), .B_i(C_s2_25_0), .c_in(C_s3_25_0), .S_o(S_s1_26_0), .c_out(C_s1_26_0));
logic S_s1_27_0, C_s1_27_0;
FA FA_s1_27_0(.A_i(S_s2_27_0), .B_i(C_s2_26_0), .c_in(C_s3_26_0), .S_o(S_s1_27_0), .c_out(C_s1_27_0));
logic S_s1_28_0, C_s1_28_0;
FA FA_s1_28_0(.A_i(S_s2_28_0), .B_i(C_s2_27_0), .c_in(C_s3_27_0), .S_o(S_s1_28_0), .c_out(C_s1_28_0));
logic S_s1_29_0, C_s1_29_0;
FA FA_s1_29_0(.A_i(S_s2_29_0), .B_i(C_s2_28_0), .c_in(C_s3_28_0), .S_o(S_s1_29_0), .c_out(C_s1_29_0));
logic S_s1_30_0, C_s1_30_0;
FA FA_s1_30_0(.A_i(S_s2_30_0), .B_i(C_s2_29_0), .c_in(C_s3_29_0), .S_o(S_s1_30_0), .c_out(C_s1_30_0));
logic S_s1_31_0, C_s1_31_0;
FA FA_s1_31_0(.A_i(S_s2_31_0), .B_i(C_s2_30_0), .c_in(C_s3_30_0), .S_o(S_s1_31_0), .c_out(C_s1_31_0));
logic S_s1_32_0, C_s1_32_0;
FA FA_s1_32_0(.A_i(S_s2_32_0), .B_i(C_s2_31_0), .c_in(C_s3_31_0), .S_o(S_s1_32_0), .c_out(C_s1_32_0));
logic S_s1_33_0, C_s1_33_0;
FA FA_s1_33_0(.A_i(S_s2_33_0), .B_i(C_s2_32_0), .c_in(C_s3_32_0), .S_o(S_s1_33_0), .c_out(C_s1_33_0));
logic S_s1_34_0, C_s1_34_0;
FA FA_s1_34_0(.A_i(S_s2_34_0), .B_i(C_s2_33_0), .c_in(C_s3_33_0), .S_o(S_s1_34_0), .c_out(C_s1_34_0));
logic S_s1_35_0, C_s1_35_0;
FA FA_s1_35_0(.A_i(S_s2_35_0), .B_i(C_s2_34_0), .c_in(C_s3_34_0), .S_o(S_s1_35_0), .c_out(C_s1_35_0));
logic S_s1_36_0, C_s1_36_0;
FA FA_s1_36_0(.A_i(S_s2_36_0), .B_i(C_s2_35_0), .c_in(C_s3_35_0), .S_o(S_s1_36_0), .c_out(C_s1_36_0));
logic S_s1_37_0, C_s1_37_0;
FA FA_s1_37_0(.A_i(S_s2_37_0), .B_i(C_s2_36_0), .c_in(C_s3_36_0), .S_o(S_s1_37_0), .c_out(C_s1_37_0));
logic S_s1_38_0, C_s1_38_0;
FA FA_s1_38_0(.A_i(S_s2_38_0), .B_i(C_s2_37_0), .c_in(C_s3_37_0), .S_o(S_s1_38_0), .c_out(C_s1_38_0));
logic S_s1_39_0, C_s1_39_0;
FA FA_s1_39_0(.A_i(S_s2_39_0), .B_i(C_s2_38_0), .c_in(C_s3_38_0), .S_o(S_s1_39_0), .c_out(C_s1_39_0));
logic S_s1_40_0, C_s1_40_0;
FA FA_s1_40_0(.A_i(S_s2_40_0), .B_i(C_s2_39_0), .c_in(C_s3_39_0), .S_o(S_s1_40_0), .c_out(C_s1_40_0));
logic S_s1_41_0, C_s1_41_0;
FA FA_s1_41_0(.A_i(S_s2_41_0), .B_i(C_s2_40_0), .c_in(C_s3_40_0), .S_o(S_s1_41_0), .c_out(C_s1_41_0));
logic S_s1_42_0, C_s1_42_0;
FA FA_s1_42_0(.A_i(S_s2_42_0), .B_i(C_s2_41_0), .c_in(C_s3_41_0), .S_o(S_s1_42_0), .c_out(C_s1_42_0));
logic S_s1_43_0, C_s1_43_0;
FA FA_s1_43_0(.A_i(S_s2_43_0), .B_i(C_s2_42_0), .c_in(C_s3_42_0), .S_o(S_s1_43_0), .c_out(C_s1_43_0));
logic S_s1_44_0, C_s1_44_0;
FA FA_s1_44_0(.A_i(S_s2_44_0), .B_i(C_s2_43_0), .c_in(C_s3_43_0), .S_o(S_s1_44_0), .c_out(C_s1_44_0));
logic S_s1_45_0, C_s1_45_0;
FA FA_s1_45_0(.A_i(S_s2_45_0), .B_i(C_s2_44_0), .c_in(C_s3_44_0), .S_o(S_s1_45_0), .c_out(C_s1_45_0));
logic S_s1_46_0, C_s1_46_0;
FA FA_s1_46_0(.A_i(S_s2_46_0), .B_i(C_s2_45_0), .c_in(C_s3_45_0), .S_o(S_s1_46_0), .c_out(C_s1_46_0));
logic S_s1_47_0, C_s1_47_0;
FA FA_s1_47_0(.A_i(S_s2_47_0), .B_i(C_s2_46_0), .c_in(C_s3_46_0), .S_o(S_s1_47_0), .c_out(C_s1_47_0));
logic S_s1_48_0, C_s1_48_0;
FA FA_s1_48_0(.A_i(S_s2_48_0), .B_i(C_s2_47_0), .c_in(C_s3_47_0), .S_o(S_s1_48_0), .c_out(C_s1_48_0));
logic S_s1_49_0, C_s1_49_0;
FA FA_s1_49_0(.A_i(S_s2_49_0), .B_i(C_s2_48_0), .c_in(C_s3_48_0), .S_o(S_s1_49_0), .c_out(C_s1_49_0));
logic S_s1_50_0, C_s1_50_0;
FA FA_s1_50_0(.A_i(S_s2_50_0), .B_i(C_s2_49_0), .c_in(C_s3_49_0), .S_o(S_s1_50_0), .c_out(C_s1_50_0));
logic S_s1_51_0, C_s1_51_0;
FA FA_s1_51_0(.A_i(S_s2_51_0), .B_i(C_s2_50_0), .c_in(C_s3_50_0), .S_o(S_s1_51_0), .c_out(C_s1_51_0));
logic S_s1_52_0, C_s1_52_0;
FA FA_s1_52_0(.A_i(S_s2_52_0), .B_i(C_s2_51_0), .c_in(C_s3_51_0), .S_o(S_s1_52_0), .c_out(C_s1_52_0));
logic S_s1_53_0, C_s1_53_0;
FA FA_s1_53_0(.A_i(S_s2_53_0), .B_i(C_s2_52_0), .c_in(C_s3_52_0), .S_o(S_s1_53_0), .c_out(C_s1_53_0));
logic S_s1_54_0, C_s1_54_0;
FA FA_s1_54_0(.A_i(S_s2_54_0), .B_i(C_s2_53_0), .c_in(C_s3_53_0), .S_o(S_s1_54_0), .c_out(C_s1_54_0));
logic S_s1_55_0, C_s1_55_0;
FA FA_s1_55_0(.A_i(S_s2_55_0), .B_i(C_s2_54_0), .c_in(C_s3_54_0), .S_o(S_s1_55_0), .c_out(C_s1_55_0));
logic S_s1_56_0, C_s1_56_0;
FA FA_s1_56_0(.A_i(S_s2_56_0), .B_i(C_s2_55_0), .c_in(C_s3_55_0), .S_o(S_s1_56_0), .c_out(C_s1_56_0));
logic S_s1_57_0, C_s1_57_0;
FA FA_s1_57_0(.A_i(S_s2_57_0), .B_i(C_s2_56_0), .c_in(C_s3_56_0), .S_o(S_s1_57_0), .c_out(C_s1_57_0));
logic S_s1_58_0, C_s1_58_0;
FA FA_s1_58_0(.A_i(S_s2_58_0), .B_i(C_s2_57_0), .c_in(C_s3_57_0), .S_o(S_s1_58_0), .c_out(C_s1_58_0));
logic S_s1_59_0, C_s1_59_0;
FA FA_s1_59_0(.A_i(S_s2_59_0), .B_i(C_s2_58_0), .c_in(comb[31][28]), .S_o(S_s1_59_0), .c_out(C_s1_59_0));
logic S_s1_60_0, C_s1_60_0;
FA FA_s1_60_0(.A_i(S_s2_60_0), .B_i(C_s2_59_0), .c_in(comb[31][29]), .S_o(S_s1_60_0), .c_out(C_s1_60_0));
logic S_s1_61_0, C_s1_61_0;
FA FA_s1_61_0(.A_i(C_s2_60_0), .B_i(comb[30][31]), .c_in(comb[31][30]), .S_o(S_s1_61_0), .c_out(C_s1_61_0));
// stage 1 end ======================================================================================================= 


// logic [63:0] last_top_row, last_bot_row;
assign row_top = {1'b0, C_s1_61_0, S_s1_61_0, S_s1_60_0, S_s1_59_0, S_s1_58_0, S_s1_57_0, S_s1_56_0, S_s1_55_0, S_s1_54_0, S_s1_53_0, S_s1_52_0, S_s1_51_0, S_s1_50_0, S_s1_49_0, S_s1_48_0, S_s1_47_0, S_s1_46_0, S_s1_45_0, S_s1_44_0, S_s1_43_0, S_s1_42_0, S_s1_41_0, S_s1_40_0, S_s1_39_0, S_s1_38_0, S_s1_37_0, S_s1_36_0, S_s1_35_0, S_s1_34_0, S_s1_33_0, S_s1_32_0, S_s1_31_0, S_s1_30_0, S_s1_29_0, S_s1_28_0, S_s1_27_0, S_s1_26_0, S_s1_25_0, S_s1_24_0, S_s1_23_0, S_s1_22_0, S_s1_21_0, S_s1_20_0, S_s1_19_0, S_s1_18_0, S_s1_17_0, S_s1_16_0, S_s1_15_0, S_s1_14_0, S_s1_13_0, S_s1_12_0, S_s1_11_0, S_s1_10_0, S_s1_9_0, S_s1_8_0, S_s1_7_0, S_s1_6_0, S_s1_5_0, S_s1_4_0, S_s1_3_0, S_s1_2_0, comb[0][1], comb[0][0]};
assign row_bot = {1'b0, comb[31][31], C_s1_60_0, C_s1_59_0, C_s1_58_0, C_s1_57_0, C_s1_56_0, C_s1_55_0, C_s1_54_0, C_s1_53_0, C_s1_52_0, C_s1_51_0, C_s1_50_0, C_s1_49_0, C_s1_48_0, C_s1_47_0, C_s1_46_0, C_s1_45_0, C_s1_44_0, C_s1_43_0, C_s1_42_0, C_s1_41_0, C_s1_40_0, C_s1_39_0, C_s1_38_0, C_s1_37_0, C_s1_36_0, C_s1_35_0, C_s1_34_0, C_s1_33_0, C_s1_32_0, C_s1_31_0, C_s1_30_0, C_s1_29_0, C_s1_28_0, C_s1_27_0, C_s1_26_0, C_s1_25_0, C_s1_24_0, C_s1_23_0, C_s1_22_0, C_s1_21_0, C_s1_20_0, C_s1_19_0, C_s1_18_0, C_s1_17_0, C_s1_16_0, C_s1_15_0, C_s1_14_0, C_s1_13_0, C_s1_12_0, C_s1_11_0, C_s1_10_0, C_s1_9_0, C_s1_8_0, C_s1_7_0, C_s1_6_0, C_s1_5_0, C_s1_4_0, C_s1_3_0, C_s1_2_0, comb[2][0], comb[1][0], 1'b0};
// assign prodAB = last_top_row + last_bot_row;    // combine and find the sum, naive implementation
endmodule
