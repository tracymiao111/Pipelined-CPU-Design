module dadda_tree(
  input logic[31:0] opA,      
  input logic[31:0] opB,      
  output logic[63:0] prodAB   
);
logic [31:0] comb[32]; 
genvar i, j; 
for(i = 0; i < 32; ++i) begin 
  for(j = 0; j < 32; ++j) begin 
      assign comb[i][j] = opA[j] & opB[i]; 
  end 
end 
logic p0000;
assign p0000 = opB[0] & opA[0];
logic p0001;
assign p0001 = opB[0] & opA[1];
logic p0002;
assign p0002 = opB[0] & opA[2];
logic p0003;
assign p0003 = opB[0] & opA[3];
logic p0004;
assign p0004 = opB[0] & opA[4];
logic p0005;
assign p0005 = opB[0] & opA[5];
logic p0006;
assign p0006 = opB[0] & opA[6];
logic p0007;
assign p0007 = opB[0] & opA[7];
logic p0008;
assign p0008 = opB[0] & opA[8];
logic p0009;
assign p0009 = opB[0] & opA[9];
logic p0010;
assign p0010 = opB[0] & opA[10];
logic p0011;
assign p0011 = opB[0] & opA[11];
logic p0012;
assign p0012 = opB[0] & opA[12];
logic p0013;
assign p0013 = opB[0] & opA[13];
logic p0014;
assign p0014 = opB[0] & opA[14];
logic p0015;
assign p0015 = opB[0] & opA[15];
logic p0016;
assign p0016 = opB[0] & opA[16];
logic p0017;
assign p0017 = opB[0] & opA[17];
logic p0018;
assign p0018 = opB[0] & opA[18];
logic p0019;
assign p0019 = opB[0] & opA[19];
logic p0020;
assign p0020 = opB[0] & opA[20];
logic p0021;
assign p0021 = opB[0] & opA[21];
logic p0022;
assign p0022 = opB[0] & opA[22];
logic p0023;
assign p0023 = opB[0] & opA[23];
logic p0024;
assign p0024 = opB[0] & opA[24];
logic p0025;
assign p0025 = opB[0] & opA[25];
logic p0026;
assign p0026 = opB[0] & opA[26];
logic p0027;
assign p0027 = opB[0] & opA[27];
logic p0028;
assign p0028 = opB[0] & opA[28];
logic p0029;
assign p0029 = opB[0] & opA[29];
logic p0030;
assign p0030 = opB[0] & opA[30];
logic p0031;
assign p0031 = opB[0] & opA[31];
logic p0100;
assign p0100 = opB[1] & opA[0];
logic p0101;
assign p0101 = opB[1] & opA[1];
logic p0102;
assign p0102 = opB[1] & opA[2];
logic p0103;
assign p0103 = opB[1] & opA[3];
logic p0104;
assign p0104 = opB[1] & opA[4];
logic p0105;
assign p0105 = opB[1] & opA[5];
logic p0106;
assign p0106 = opB[1] & opA[6];
logic p0107;
assign p0107 = opB[1] & opA[7];
logic p0108;
assign p0108 = opB[1] & opA[8];
logic p0109;
assign p0109 = opB[1] & opA[9];
logic p0110;
assign p0110 = opB[1] & opA[10];
logic p0111;
assign p0111 = opB[1] & opA[11];
logic p0112;
assign p0112 = opB[1] & opA[12];
logic p0113;
assign p0113 = opB[1] & opA[13];
logic p0114;
assign p0114 = opB[1] & opA[14];
logic p0115;
assign p0115 = opB[1] & opA[15];
logic p0116;
assign p0116 = opB[1] & opA[16];
logic p0117;
assign p0117 = opB[1] & opA[17];
logic p0118;
assign p0118 = opB[1] & opA[18];
logic p0119;
assign p0119 = opB[1] & opA[19];
logic p0120;
assign p0120 = opB[1] & opA[20];
logic p0121;
assign p0121 = opB[1] & opA[21];
logic p0122;
assign p0122 = opB[1] & opA[22];
logic p0123;
assign p0123 = opB[1] & opA[23];
logic p0124;
assign p0124 = opB[1] & opA[24];
logic p0125;
assign p0125 = opB[1] & opA[25];
logic p0126;
assign p0126 = opB[1] & opA[26];
logic p0127;
assign p0127 = opB[1] & opA[27];
logic p0128;
assign p0128 = opB[1] & opA[28];
logic p0129;
assign p0129 = opB[1] & opA[29];
logic p0130;
assign p0130 = opB[1] & opA[30];
logic p0131;
assign p0131 = opB[1] & opA[31];
logic p0200;
assign p0200 = opB[2] & opA[0];
logic p0201;
assign p0201 = opB[2] & opA[1];
logic p0202;
assign p0202 = opB[2] & opA[2];
logic p0203;
assign p0203 = opB[2] & opA[3];
logic p0204;
assign p0204 = opB[2] & opA[4];
logic p0205;
assign p0205 = opB[2] & opA[5];
logic p0206;
assign p0206 = opB[2] & opA[6];
logic p0207;
assign p0207 = opB[2] & opA[7];
logic p0208;
assign p0208 = opB[2] & opA[8];
logic p0209;
assign p0209 = opB[2] & opA[9];
logic p0210;
assign p0210 = opB[2] & opA[10];
logic p0211;
assign p0211 = opB[2] & opA[11];
logic p0212;
assign p0212 = opB[2] & opA[12];
logic p0213;
assign p0213 = opB[2] & opA[13];
logic p0214;
assign p0214 = opB[2] & opA[14];
logic p0215;
assign p0215 = opB[2] & opA[15];
logic p0216;
assign p0216 = opB[2] & opA[16];
logic p0217;
assign p0217 = opB[2] & opA[17];
logic p0218;
assign p0218 = opB[2] & opA[18];
logic p0219;
assign p0219 = opB[2] & opA[19];
logic p0220;
assign p0220 = opB[2] & opA[20];
logic p0221;
assign p0221 = opB[2] & opA[21];
logic p0222;
assign p0222 = opB[2] & opA[22];
logic p0223;
assign p0223 = opB[2] & opA[23];
logic p0224;
assign p0224 = opB[2] & opA[24];
logic p0225;
assign p0225 = opB[2] & opA[25];
logic p0226;
assign p0226 = opB[2] & opA[26];
logic p0227;
assign p0227 = opB[2] & opA[27];
logic p0228;
assign p0228 = opB[2] & opA[28];
logic p0229;
assign p0229 = opB[2] & opA[29];
logic p0230;
assign p0230 = opB[2] & opA[30];
logic p0231;
assign p0231 = opB[2] & opA[31];
logic p0300;
assign p0300 = opB[3] & opA[0];
logic p0301;
assign p0301 = opB[3] & opA[1];
logic p0302;
assign p0302 = opB[3] & opA[2];
logic p0303;
assign p0303 = opB[3] & opA[3];
logic p0304;
assign p0304 = opB[3] & opA[4];
logic p0305;
assign p0305 = opB[3] & opA[5];
logic p0306;
assign p0306 = opB[3] & opA[6];
logic p0307;
assign p0307 = opB[3] & opA[7];
logic p0308;
assign p0308 = opB[3] & opA[8];
logic p0309;
assign p0309 = opB[3] & opA[9];
logic p0310;
assign p0310 = opB[3] & opA[10];
logic p0311;
assign p0311 = opB[3] & opA[11];
logic p0312;
assign p0312 = opB[3] & opA[12];
logic p0313;
assign p0313 = opB[3] & opA[13];
logic p0314;
assign p0314 = opB[3] & opA[14];
logic p0315;
assign p0315 = opB[3] & opA[15];
logic p0316;
assign p0316 = opB[3] & opA[16];
logic p0317;
assign p0317 = opB[3] & opA[17];
logic p0318;
assign p0318 = opB[3] & opA[18];
logic p0319;
assign p0319 = opB[3] & opA[19];
logic p0320;
assign p0320 = opB[3] & opA[20];
logic p0321;
assign p0321 = opB[3] & opA[21];
logic p0322;
assign p0322 = opB[3] & opA[22];
logic p0323;
assign p0323 = opB[3] & opA[23];
logic p0324;
assign p0324 = opB[3] & opA[24];
logic p0325;
assign p0325 = opB[3] & opA[25];
logic p0326;
assign p0326 = opB[3] & opA[26];
logic p0327;
assign p0327 = opB[3] & opA[27];
logic p0328;
assign p0328 = opB[3] & opA[28];
logic p0329;
assign p0329 = opB[3] & opA[29];
logic p0330;
assign p0330 = opB[3] & opA[30];
logic p0331;
assign p0331 = opB[3] & opA[31];
logic p0400;
assign p0400 = opB[4] & opA[0];
logic p0401;
assign p0401 = opB[4] & opA[1];
logic p0402;
assign p0402 = opB[4] & opA[2];
logic p0403;
assign p0403 = opB[4] & opA[3];
logic p0404;
assign p0404 = opB[4] & opA[4];
logic p0405;
assign p0405 = opB[4] & opA[5];
logic p0406;
assign p0406 = opB[4] & opA[6];
logic p0407;
assign p0407 = opB[4] & opA[7];
logic p0408;
assign p0408 = opB[4] & opA[8];
logic p0409;
assign p0409 = opB[4] & opA[9];
logic p0410;
assign p0410 = opB[4] & opA[10];
logic p0411;
assign p0411 = opB[4] & opA[11];
logic p0412;
assign p0412 = opB[4] & opA[12];
logic p0413;
assign p0413 = opB[4] & opA[13];
logic p0414;
assign p0414 = opB[4] & opA[14];
logic p0415;
assign p0415 = opB[4] & opA[15];
logic p0416;
assign p0416 = opB[4] & opA[16];
logic p0417;
assign p0417 = opB[4] & opA[17];
logic p0418;
assign p0418 = opB[4] & opA[18];
logic p0419;
assign p0419 = opB[4] & opA[19];
logic p0420;
assign p0420 = opB[4] & opA[20];
logic p0421;
assign p0421 = opB[4] & opA[21];
logic p0422;
assign p0422 = opB[4] & opA[22];
logic p0423;
assign p0423 = opB[4] & opA[23];
logic p0424;
assign p0424 = opB[4] & opA[24];
logic p0425;
assign p0425 = opB[4] & opA[25];
logic p0426;
assign p0426 = opB[4] & opA[26];
logic p0427;
assign p0427 = opB[4] & opA[27];
logic p0428;
assign p0428 = opB[4] & opA[28];
logic p0429;
assign p0429 = opB[4] & opA[29];
logic p0430;
assign p0430 = opB[4] & opA[30];
logic p0431;
assign p0431 = opB[4] & opA[31];
logic p0500;
assign p0500 = opB[5] & opA[0];
logic p0501;
assign p0501 = opB[5] & opA[1];
logic p0502;
assign p0502 = opB[5] & opA[2];
logic p0503;
assign p0503 = opB[5] & opA[3];
logic p0504;
assign p0504 = opB[5] & opA[4];
logic p0505;
assign p0505 = opB[5] & opA[5];
logic p0506;
assign p0506 = opB[5] & opA[6];
logic p0507;
assign p0507 = opB[5] & opA[7];
logic p0508;
assign p0508 = opB[5] & opA[8];
logic p0509;
assign p0509 = opB[5] & opA[9];
logic p0510;
assign p0510 = opB[5] & opA[10];
logic p0511;
assign p0511 = opB[5] & opA[11];
logic p0512;
assign p0512 = opB[5] & opA[12];
logic p0513;
assign p0513 = opB[5] & opA[13];
logic p0514;
assign p0514 = opB[5] & opA[14];
logic p0515;
assign p0515 = opB[5] & opA[15];
logic p0516;
assign p0516 = opB[5] & opA[16];
logic p0517;
assign p0517 = opB[5] & opA[17];
logic p0518;
assign p0518 = opB[5] & opA[18];
logic p0519;
assign p0519 = opB[5] & opA[19];
logic p0520;
assign p0520 = opB[5] & opA[20];
logic p0521;
assign p0521 = opB[5] & opA[21];
logic p0522;
assign p0522 = opB[5] & opA[22];
logic p0523;
assign p0523 = opB[5] & opA[23];
logic p0524;
assign p0524 = opB[5] & opA[24];
logic p0525;
assign p0525 = opB[5] & opA[25];
logic p0526;
assign p0526 = opB[5] & opA[26];
logic p0527;
assign p0527 = opB[5] & opA[27];
logic p0528;
assign p0528 = opB[5] & opA[28];
logic p0529;
assign p0529 = opB[5] & opA[29];
logic p0530;
assign p0530 = opB[5] & opA[30];
logic p0531;
assign p0531 = opB[5] & opA[31];
logic p0600;
assign p0600 = opB[6] & opA[0];
logic p0601;
assign p0601 = opB[6] & opA[1];
logic p0602;
assign p0602 = opB[6] & opA[2];
logic p0603;
assign p0603 = opB[6] & opA[3];
logic p0604;
assign p0604 = opB[6] & opA[4];
logic p0605;
assign p0605 = opB[6] & opA[5];
logic p0606;
assign p0606 = opB[6] & opA[6];
logic p0607;
assign p0607 = opB[6] & opA[7];
logic p0608;
assign p0608 = opB[6] & opA[8];
logic p0609;
assign p0609 = opB[6] & opA[9];
logic p0610;
assign p0610 = opB[6] & opA[10];
logic p0611;
assign p0611 = opB[6] & opA[11];
logic p0612;
assign p0612 = opB[6] & opA[12];
logic p0613;
assign p0613 = opB[6] & opA[13];
logic p0614;
assign p0614 = opB[6] & opA[14];
logic p0615;
assign p0615 = opB[6] & opA[15];
logic p0616;
assign p0616 = opB[6] & opA[16];
logic p0617;
assign p0617 = opB[6] & opA[17];
logic p0618;
assign p0618 = opB[6] & opA[18];
logic p0619;
assign p0619 = opB[6] & opA[19];
logic p0620;
assign p0620 = opB[6] & opA[20];
logic p0621;
assign p0621 = opB[6] & opA[21];
logic p0622;
assign p0622 = opB[6] & opA[22];
logic p0623;
assign p0623 = opB[6] & opA[23];
logic p0624;
assign p0624 = opB[6] & opA[24];
logic p0625;
assign p0625 = opB[6] & opA[25];
logic p0626;
assign p0626 = opB[6] & opA[26];
logic p0627;
assign p0627 = opB[6] & opA[27];
logic p0628;
assign p0628 = opB[6] & opA[28];
logic p0629;
assign p0629 = opB[6] & opA[29];
logic p0630;
assign p0630 = opB[6] & opA[30];
logic p0631;
assign p0631 = opB[6] & opA[31];
logic p0700;
assign p0700 = opB[7] & opA[0];
logic p0701;
assign p0701 = opB[7] & opA[1];
logic p0702;
assign p0702 = opB[7] & opA[2];
logic p0703;
assign p0703 = opB[7] & opA[3];
logic p0704;
assign p0704 = opB[7] & opA[4];
logic p0705;
assign p0705 = opB[7] & opA[5];
logic p0706;
assign p0706 = opB[7] & opA[6];
logic p0707;
assign p0707 = opB[7] & opA[7];
logic p0708;
assign p0708 = opB[7] & opA[8];
logic p0709;
assign p0709 = opB[7] & opA[9];
logic p0710;
assign p0710 = opB[7] & opA[10];
logic p0711;
assign p0711 = opB[7] & opA[11];
logic p0712;
assign p0712 = opB[7] & opA[12];
logic p0713;
assign p0713 = opB[7] & opA[13];
logic p0714;
assign p0714 = opB[7] & opA[14];
logic p0715;
assign p0715 = opB[7] & opA[15];
logic p0716;
assign p0716 = opB[7] & opA[16];
logic p0717;
assign p0717 = opB[7] & opA[17];
logic p0718;
assign p0718 = opB[7] & opA[18];
logic p0719;
assign p0719 = opB[7] & opA[19];
logic p0720;
assign p0720 = opB[7] & opA[20];
logic p0721;
assign p0721 = opB[7] & opA[21];
logic p0722;
assign p0722 = opB[7] & opA[22];
logic p0723;
assign p0723 = opB[7] & opA[23];
logic p0724;
assign p0724 = opB[7] & opA[24];
logic p0725;
assign p0725 = opB[7] & opA[25];
logic p0726;
assign p0726 = opB[7] & opA[26];
logic p0727;
assign p0727 = opB[7] & opA[27];
logic p0728;
assign p0728 = opB[7] & opA[28];
logic p0729;
assign p0729 = opB[7] & opA[29];
logic p0730;
assign p0730 = opB[7] & opA[30];
logic p0731;
assign p0731 = opB[7] & opA[31];
logic p0800;
assign p0800 = opB[8] & opA[0];
logic p0801;
assign p0801 = opB[8] & opA[1];
logic p0802;
assign p0802 = opB[8] & opA[2];
logic p0803;
assign p0803 = opB[8] & opA[3];
logic p0804;
assign p0804 = opB[8] & opA[4];
logic p0805;
assign p0805 = opB[8] & opA[5];
logic p0806;
assign p0806 = opB[8] & opA[6];
logic p0807;
assign p0807 = opB[8] & opA[7];
logic p0808;
assign p0808 = opB[8] & opA[8];
logic p0809;
assign p0809 = opB[8] & opA[9];
logic p0810;
assign p0810 = opB[8] & opA[10];
logic p0811;
assign p0811 = opB[8] & opA[11];
logic p0812;
assign p0812 = opB[8] & opA[12];
logic p0813;
assign p0813 = opB[8] & opA[13];
logic p0814;
assign p0814 = opB[8] & opA[14];
logic p0815;
assign p0815 = opB[8] & opA[15];
logic p0816;
assign p0816 = opB[8] & opA[16];
logic p0817;
assign p0817 = opB[8] & opA[17];
logic p0818;
assign p0818 = opB[8] & opA[18];
logic p0819;
assign p0819 = opB[8] & opA[19];
logic p0820;
assign p0820 = opB[8] & opA[20];
logic p0821;
assign p0821 = opB[8] & opA[21];
logic p0822;
assign p0822 = opB[8] & opA[22];
logic p0823;
assign p0823 = opB[8] & opA[23];
logic p0824;
assign p0824 = opB[8] & opA[24];
logic p0825;
assign p0825 = opB[8] & opA[25];
logic p0826;
assign p0826 = opB[8] & opA[26];
logic p0827;
assign p0827 = opB[8] & opA[27];
logic p0828;
assign p0828 = opB[8] & opA[28];
logic p0829;
assign p0829 = opB[8] & opA[29];
logic p0830;
assign p0830 = opB[8] & opA[30];
logic p0831;
assign p0831 = opB[8] & opA[31];
logic p0900;
assign p0900 = opB[9] & opA[0];
logic p0901;
assign p0901 = opB[9] & opA[1];
logic p0902;
assign p0902 = opB[9] & opA[2];
logic p0903;
assign p0903 = opB[9] & opA[3];
logic p0904;
assign p0904 = opB[9] & opA[4];
logic p0905;
assign p0905 = opB[9] & opA[5];
logic p0906;
assign p0906 = opB[9] & opA[6];
logic p0907;
assign p0907 = opB[9] & opA[7];
logic p0908;
assign p0908 = opB[9] & opA[8];
logic p0909;
assign p0909 = opB[9] & opA[9];
logic p0910;
assign p0910 = opB[9] & opA[10];
logic p0911;
assign p0911 = opB[9] & opA[11];
logic p0912;
assign p0912 = opB[9] & opA[12];
logic p0913;
assign p0913 = opB[9] & opA[13];
logic p0914;
assign p0914 = opB[9] & opA[14];
logic p0915;
assign p0915 = opB[9] & opA[15];
logic p0916;
assign p0916 = opB[9] & opA[16];
logic p0917;
assign p0917 = opB[9] & opA[17];
logic p0918;
assign p0918 = opB[9] & opA[18];
logic p0919;
assign p0919 = opB[9] & opA[19];
logic p0920;
assign p0920 = opB[9] & opA[20];
logic p0921;
assign p0921 = opB[9] & opA[21];
logic p0922;
assign p0922 = opB[9] & opA[22];
logic p0923;
assign p0923 = opB[9] & opA[23];
logic p0924;
assign p0924 = opB[9] & opA[24];
logic p0925;
assign p0925 = opB[9] & opA[25];
logic p0926;
assign p0926 = opB[9] & opA[26];
logic p0927;
assign p0927 = opB[9] & opA[27];
logic p0928;
assign p0928 = opB[9] & opA[28];
logic p0929;
assign p0929 = opB[9] & opA[29];
logic p0930;
assign p0930 = opB[9] & opA[30];
logic p0931;
assign p0931 = opB[9] & opA[31];
logic p1000;
assign p1000 = opB[10] & opA[0];
logic p1001;
assign p1001 = opB[10] & opA[1];
logic p1002;
assign p1002 = opB[10] & opA[2];
logic p1003;
assign p1003 = opB[10] & opA[3];
logic p1004;
assign p1004 = opB[10] & opA[4];
logic p1005;
assign p1005 = opB[10] & opA[5];
logic p1006;
assign p1006 = opB[10] & opA[6];
logic p1007;
assign p1007 = opB[10] & opA[7];
logic p1008;
assign p1008 = opB[10] & opA[8];
logic p1009;
assign p1009 = opB[10] & opA[9];
logic p1010;
assign p1010 = opB[10] & opA[10];
logic p1011;
assign p1011 = opB[10] & opA[11];
logic p1012;
assign p1012 = opB[10] & opA[12];
logic p1013;
assign p1013 = opB[10] & opA[13];
logic p1014;
assign p1014 = opB[10] & opA[14];
logic p1015;
assign p1015 = opB[10] & opA[15];
logic p1016;
assign p1016 = opB[10] & opA[16];
logic p1017;
assign p1017 = opB[10] & opA[17];
logic p1018;
assign p1018 = opB[10] & opA[18];
logic p1019;
assign p1019 = opB[10] & opA[19];
logic p1020;
assign p1020 = opB[10] & opA[20];
logic p1021;
assign p1021 = opB[10] & opA[21];
logic p1022;
assign p1022 = opB[10] & opA[22];
logic p1023;
assign p1023 = opB[10] & opA[23];
logic p1024;
assign p1024 = opB[10] & opA[24];
logic p1025;
assign p1025 = opB[10] & opA[25];
logic p1026;
assign p1026 = opB[10] & opA[26];
logic p1027;
assign p1027 = opB[10] & opA[27];
logic p1028;
assign p1028 = opB[10] & opA[28];
logic p1029;
assign p1029 = opB[10] & opA[29];
logic p1030;
assign p1030 = opB[10] & opA[30];
logic p1031;
assign p1031 = opB[10] & opA[31];
logic p1100;
assign p1100 = opB[11] & opA[0];
logic p1101;
assign p1101 = opB[11] & opA[1];
logic p1102;
assign p1102 = opB[11] & opA[2];
logic p1103;
assign p1103 = opB[11] & opA[3];
logic p1104;
assign p1104 = opB[11] & opA[4];
logic p1105;
assign p1105 = opB[11] & opA[5];
logic p1106;
assign p1106 = opB[11] & opA[6];
logic p1107;
assign p1107 = opB[11] & opA[7];
logic p1108;
assign p1108 = opB[11] & opA[8];
logic p1109;
assign p1109 = opB[11] & opA[9];
logic p1110;
assign p1110 = opB[11] & opA[10];
logic p1111;
assign p1111 = opB[11] & opA[11];
logic p1112;
assign p1112 = opB[11] & opA[12];
logic p1113;
assign p1113 = opB[11] & opA[13];
logic p1114;
assign p1114 = opB[11] & opA[14];
logic p1115;
assign p1115 = opB[11] & opA[15];
logic p1116;
assign p1116 = opB[11] & opA[16];
logic p1117;
assign p1117 = opB[11] & opA[17];
logic p1118;
assign p1118 = opB[11] & opA[18];
logic p1119;
assign p1119 = opB[11] & opA[19];
logic p1120;
assign p1120 = opB[11] & opA[20];
logic p1121;
assign p1121 = opB[11] & opA[21];
logic p1122;
assign p1122 = opB[11] & opA[22];
logic p1123;
assign p1123 = opB[11] & opA[23];
logic p1124;
assign p1124 = opB[11] & opA[24];
logic p1125;
assign p1125 = opB[11] & opA[25];
logic p1126;
assign p1126 = opB[11] & opA[26];
logic p1127;
assign p1127 = opB[11] & opA[27];
logic p1128;
assign p1128 = opB[11] & opA[28];
logic p1129;
assign p1129 = opB[11] & opA[29];
logic p1130;
assign p1130 = opB[11] & opA[30];
logic p1131;
assign p1131 = opB[11] & opA[31];
logic p1200;
assign p1200 = opB[12] & opA[0];
logic p1201;
assign p1201 = opB[12] & opA[1];
logic p1202;
assign p1202 = opB[12] & opA[2];
logic p1203;
assign p1203 = opB[12] & opA[3];
logic p1204;
assign p1204 = opB[12] & opA[4];
logic p1205;
assign p1205 = opB[12] & opA[5];
logic p1206;
assign p1206 = opB[12] & opA[6];
logic p1207;
assign p1207 = opB[12] & opA[7];
logic p1208;
assign p1208 = opB[12] & opA[8];
logic p1209;
assign p1209 = opB[12] & opA[9];
logic p1210;
assign p1210 = opB[12] & opA[10];
logic p1211;
assign p1211 = opB[12] & opA[11];
logic p1212;
assign p1212 = opB[12] & opA[12];
logic p1213;
assign p1213 = opB[12] & opA[13];
logic p1214;
assign p1214 = opB[12] & opA[14];
logic p1215;
assign p1215 = opB[12] & opA[15];
logic p1216;
assign p1216 = opB[12] & opA[16];
logic p1217;
assign p1217 = opB[12] & opA[17];
logic p1218;
assign p1218 = opB[12] & opA[18];
logic p1219;
assign p1219 = opB[12] & opA[19];
logic p1220;
assign p1220 = opB[12] & opA[20];
logic p1221;
assign p1221 = opB[12] & opA[21];
logic p1222;
assign p1222 = opB[12] & opA[22];
logic p1223;
assign p1223 = opB[12] & opA[23];
logic p1224;
assign p1224 = opB[12] & opA[24];
logic p1225;
assign p1225 = opB[12] & opA[25];
logic p1226;
assign p1226 = opB[12] & opA[26];
logic p1227;
assign p1227 = opB[12] & opA[27];
logic p1228;
assign p1228 = opB[12] & opA[28];
logic p1229;
assign p1229 = opB[12] & opA[29];
logic p1230;
assign p1230 = opB[12] & opA[30];
logic p1231;
assign p1231 = opB[12] & opA[31];
logic p1300;
assign p1300 = opB[13] & opA[0];
logic p1301;
assign p1301 = opB[13] & opA[1];
logic p1302;
assign p1302 = opB[13] & opA[2];
logic p1303;
assign p1303 = opB[13] & opA[3];
logic p1304;
assign p1304 = opB[13] & opA[4];
logic p1305;
assign p1305 = opB[13] & opA[5];
logic p1306;
assign p1306 = opB[13] & opA[6];
logic p1307;
assign p1307 = opB[13] & opA[7];
logic p1308;
assign p1308 = opB[13] & opA[8];
logic p1309;
assign p1309 = opB[13] & opA[9];
logic p1310;
assign p1310 = opB[13] & opA[10];
logic p1311;
assign p1311 = opB[13] & opA[11];
logic p1312;
assign p1312 = opB[13] & opA[12];
logic p1313;
assign p1313 = opB[13] & opA[13];
logic p1314;
assign p1314 = opB[13] & opA[14];
logic p1315;
assign p1315 = opB[13] & opA[15];
logic p1316;
assign p1316 = opB[13] & opA[16];
logic p1317;
assign p1317 = opB[13] & opA[17];
logic p1318;
assign p1318 = opB[13] & opA[18];
logic p1319;
assign p1319 = opB[13] & opA[19];
logic p1320;
assign p1320 = opB[13] & opA[20];
logic p1321;
assign p1321 = opB[13] & opA[21];
logic p1322;
assign p1322 = opB[13] & opA[22];
logic p1323;
assign p1323 = opB[13] & opA[23];
logic p1324;
assign p1324 = opB[13] & opA[24];
logic p1325;
assign p1325 = opB[13] & opA[25];
logic p1326;
assign p1326 = opB[13] & opA[26];
logic p1327;
assign p1327 = opB[13] & opA[27];
logic p1328;
assign p1328 = opB[13] & opA[28];
logic p1329;
assign p1329 = opB[13] & opA[29];
logic p1330;
assign p1330 = opB[13] & opA[30];
logic p1331;
assign p1331 = opB[13] & opA[31];
logic p1400;
assign p1400 = opB[14] & opA[0];
logic p1401;
assign p1401 = opB[14] & opA[1];
logic p1402;
assign p1402 = opB[14] & opA[2];
logic p1403;
assign p1403 = opB[14] & opA[3];
logic p1404;
assign p1404 = opB[14] & opA[4];
logic p1405;
assign p1405 = opB[14] & opA[5];
logic p1406;
assign p1406 = opB[14] & opA[6];
logic p1407;
assign p1407 = opB[14] & opA[7];
logic p1408;
assign p1408 = opB[14] & opA[8];
logic p1409;
assign p1409 = opB[14] & opA[9];
logic p1410;
assign p1410 = opB[14] & opA[10];
logic p1411;
assign p1411 = opB[14] & opA[11];
logic p1412;
assign p1412 = opB[14] & opA[12];
logic p1413;
assign p1413 = opB[14] & opA[13];
logic p1414;
assign p1414 = opB[14] & opA[14];
logic p1415;
assign p1415 = opB[14] & opA[15];
logic p1416;
assign p1416 = opB[14] & opA[16];
logic p1417;
assign p1417 = opB[14] & opA[17];
logic p1418;
assign p1418 = opB[14] & opA[18];
logic p1419;
assign p1419 = opB[14] & opA[19];
logic p1420;
assign p1420 = opB[14] & opA[20];
logic p1421;
assign p1421 = opB[14] & opA[21];
logic p1422;
assign p1422 = opB[14] & opA[22];
logic p1423;
assign p1423 = opB[14] & opA[23];
logic p1424;
assign p1424 = opB[14] & opA[24];
logic p1425;
assign p1425 = opB[14] & opA[25];
logic p1426;
assign p1426 = opB[14] & opA[26];
logic p1427;
assign p1427 = opB[14] & opA[27];
logic p1428;
assign p1428 = opB[14] & opA[28];
logic p1429;
assign p1429 = opB[14] & opA[29];
logic p1430;
assign p1430 = opB[14] & opA[30];
logic p1431;
assign p1431 = opB[14] & opA[31];
logic p1500;
assign p1500 = opB[15] & opA[0];
logic p1501;
assign p1501 = opB[15] & opA[1];
logic p1502;
assign p1502 = opB[15] & opA[2];
logic p1503;
assign p1503 = opB[15] & opA[3];
logic p1504;
assign p1504 = opB[15] & opA[4];
logic p1505;
assign p1505 = opB[15] & opA[5];
logic p1506;
assign p1506 = opB[15] & opA[6];
logic p1507;
assign p1507 = opB[15] & opA[7];
logic p1508;
assign p1508 = opB[15] & opA[8];
logic p1509;
assign p1509 = opB[15] & opA[9];
logic p1510;
assign p1510 = opB[15] & opA[10];
logic p1511;
assign p1511 = opB[15] & opA[11];
logic p1512;
assign p1512 = opB[15] & opA[12];
logic p1513;
assign p1513 = opB[15] & opA[13];
logic p1514;
assign p1514 = opB[15] & opA[14];
logic p1515;
assign p1515 = opB[15] & opA[15];
logic p1516;
assign p1516 = opB[15] & opA[16];
logic p1517;
assign p1517 = opB[15] & opA[17];
logic p1518;
assign p1518 = opB[15] & opA[18];
logic p1519;
assign p1519 = opB[15] & opA[19];
logic p1520;
assign p1520 = opB[15] & opA[20];
logic p1521;
assign p1521 = opB[15] & opA[21];
logic p1522;
assign p1522 = opB[15] & opA[22];
logic p1523;
assign p1523 = opB[15] & opA[23];
logic p1524;
assign p1524 = opB[15] & opA[24];
logic p1525;
assign p1525 = opB[15] & opA[25];
logic p1526;
assign p1526 = opB[15] & opA[26];
logic p1527;
assign p1527 = opB[15] & opA[27];
logic p1528;
assign p1528 = opB[15] & opA[28];
logic p1529;
assign p1529 = opB[15] & opA[29];
logic p1530;
assign p1530 = opB[15] & opA[30];
logic p1531;
assign p1531 = opB[15] & opA[31];
logic p1600;
assign p1600 = opB[16] & opA[0];
logic p1601;
assign p1601 = opB[16] & opA[1];
logic p1602;
assign p1602 = opB[16] & opA[2];
logic p1603;
assign p1603 = opB[16] & opA[3];
logic p1604;
assign p1604 = opB[16] & opA[4];
logic p1605;
assign p1605 = opB[16] & opA[5];
logic p1606;
assign p1606 = opB[16] & opA[6];
logic p1607;
assign p1607 = opB[16] & opA[7];
logic p1608;
assign p1608 = opB[16] & opA[8];
logic p1609;
assign p1609 = opB[16] & opA[9];
logic p1610;
assign p1610 = opB[16] & opA[10];
logic p1611;
assign p1611 = opB[16] & opA[11];
logic p1612;
assign p1612 = opB[16] & opA[12];
logic p1613;
assign p1613 = opB[16] & opA[13];
logic p1614;
assign p1614 = opB[16] & opA[14];
logic p1615;
assign p1615 = opB[16] & opA[15];
logic p1616;
assign p1616 = opB[16] & opA[16];
logic p1617;
assign p1617 = opB[16] & opA[17];
logic p1618;
assign p1618 = opB[16] & opA[18];
logic p1619;
assign p1619 = opB[16] & opA[19];
logic p1620;
assign p1620 = opB[16] & opA[20];
logic p1621;
assign p1621 = opB[16] & opA[21];
logic p1622;
assign p1622 = opB[16] & opA[22];
logic p1623;
assign p1623 = opB[16] & opA[23];
logic p1624;
assign p1624 = opB[16] & opA[24];
logic p1625;
assign p1625 = opB[16] & opA[25];
logic p1626;
assign p1626 = opB[16] & opA[26];
logic p1627;
assign p1627 = opB[16] & opA[27];
logic p1628;
assign p1628 = opB[16] & opA[28];
logic p1629;
assign p1629 = opB[16] & opA[29];
logic p1630;
assign p1630 = opB[16] & opA[30];
logic p1631;
assign p1631 = opB[16] & opA[31];
logic p1700;
assign p1700 = opB[17] & opA[0];
logic p1701;
assign p1701 = opB[17] & opA[1];
logic p1702;
assign p1702 = opB[17] & opA[2];
logic p1703;
assign p1703 = opB[17] & opA[3];
logic p1704;
assign p1704 = opB[17] & opA[4];
logic p1705;
assign p1705 = opB[17] & opA[5];
logic p1706;
assign p1706 = opB[17] & opA[6];
logic p1707;
assign p1707 = opB[17] & opA[7];
logic p1708;
assign p1708 = opB[17] & opA[8];
logic p1709;
assign p1709 = opB[17] & opA[9];
logic p1710;
assign p1710 = opB[17] & opA[10];
logic p1711;
assign p1711 = opB[17] & opA[11];
logic p1712;
assign p1712 = opB[17] & opA[12];
logic p1713;
assign p1713 = opB[17] & opA[13];
logic p1714;
assign p1714 = opB[17] & opA[14];
logic p1715;
assign p1715 = opB[17] & opA[15];
logic p1716;
assign p1716 = opB[17] & opA[16];
logic p1717;
assign p1717 = opB[17] & opA[17];
logic p1718;
assign p1718 = opB[17] & opA[18];
logic p1719;
assign p1719 = opB[17] & opA[19];
logic p1720;
assign p1720 = opB[17] & opA[20];
logic p1721;
assign p1721 = opB[17] & opA[21];
logic p1722;
assign p1722 = opB[17] & opA[22];
logic p1723;
assign p1723 = opB[17] & opA[23];
logic p1724;
assign p1724 = opB[17] & opA[24];
logic p1725;
assign p1725 = opB[17] & opA[25];
logic p1726;
assign p1726 = opB[17] & opA[26];
logic p1727;
assign p1727 = opB[17] & opA[27];
logic p1728;
assign p1728 = opB[17] & opA[28];
logic p1729;
assign p1729 = opB[17] & opA[29];
logic p1730;
assign p1730 = opB[17] & opA[30];
logic p1731;
assign p1731 = opB[17] & opA[31];
logic p1800;
assign p1800 = opB[18] & opA[0];
logic p1801;
assign p1801 = opB[18] & opA[1];
logic p1802;
assign p1802 = opB[18] & opA[2];
logic p1803;
assign p1803 = opB[18] & opA[3];
logic p1804;
assign p1804 = opB[18] & opA[4];
logic p1805;
assign p1805 = opB[18] & opA[5];
logic p1806;
assign p1806 = opB[18] & opA[6];
logic p1807;
assign p1807 = opB[18] & opA[7];
logic p1808;
assign p1808 = opB[18] & opA[8];
logic p1809;
assign p1809 = opB[18] & opA[9];
logic p1810;
assign p1810 = opB[18] & opA[10];
logic p1811;
assign p1811 = opB[18] & opA[11];
logic p1812;
assign p1812 = opB[18] & opA[12];
logic p1813;
assign p1813 = opB[18] & opA[13];
logic p1814;
assign p1814 = opB[18] & opA[14];
logic p1815;
assign p1815 = opB[18] & opA[15];
logic p1816;
assign p1816 = opB[18] & opA[16];
logic p1817;
assign p1817 = opB[18] & opA[17];
logic p1818;
assign p1818 = opB[18] & opA[18];
logic p1819;
assign p1819 = opB[18] & opA[19];
logic p1820;
assign p1820 = opB[18] & opA[20];
logic p1821;
assign p1821 = opB[18] & opA[21];
logic p1822;
assign p1822 = opB[18] & opA[22];
logic p1823;
assign p1823 = opB[18] & opA[23];
logic p1824;
assign p1824 = opB[18] & opA[24];
logic p1825;
assign p1825 = opB[18] & opA[25];
logic p1826;
assign p1826 = opB[18] & opA[26];
logic p1827;
assign p1827 = opB[18] & opA[27];
logic p1828;
assign p1828 = opB[18] & opA[28];
logic p1829;
assign p1829 = opB[18] & opA[29];
logic p1830;
assign p1830 = opB[18] & opA[30];
logic p1831;
assign p1831 = opB[18] & opA[31];
logic p1900;
assign p1900 = opB[19] & opA[0];
logic p1901;
assign p1901 = opB[19] & opA[1];
logic p1902;
assign p1902 = opB[19] & opA[2];
logic p1903;
assign p1903 = opB[19] & opA[3];
logic p1904;
assign p1904 = opB[19] & opA[4];
logic p1905;
assign p1905 = opB[19] & opA[5];
logic p1906;
assign p1906 = opB[19] & opA[6];
logic p1907;
assign p1907 = opB[19] & opA[7];
logic p1908;
assign p1908 = opB[19] & opA[8];
logic p1909;
assign p1909 = opB[19] & opA[9];
logic p1910;
assign p1910 = opB[19] & opA[10];
logic p1911;
assign p1911 = opB[19] & opA[11];
logic p1912;
assign p1912 = opB[19] & opA[12];
logic p1913;
assign p1913 = opB[19] & opA[13];
logic p1914;
assign p1914 = opB[19] & opA[14];
logic p1915;
assign p1915 = opB[19] & opA[15];
logic p1916;
assign p1916 = opB[19] & opA[16];
logic p1917;
assign p1917 = opB[19] & opA[17];
logic p1918;
assign p1918 = opB[19] & opA[18];
logic p1919;
assign p1919 = opB[19] & opA[19];
logic p1920;
assign p1920 = opB[19] & opA[20];
logic p1921;
assign p1921 = opB[19] & opA[21];
logic p1922;
assign p1922 = opB[19] & opA[22];
logic p1923;
assign p1923 = opB[19] & opA[23];
logic p1924;
assign p1924 = opB[19] & opA[24];
logic p1925;
assign p1925 = opB[19] & opA[25];
logic p1926;
assign p1926 = opB[19] & opA[26];
logic p1927;
assign p1927 = opB[19] & opA[27];
logic p1928;
assign p1928 = opB[19] & opA[28];
logic p1929;
assign p1929 = opB[19] & opA[29];
logic p1930;
assign p1930 = opB[19] & opA[30];
logic p1931;
assign p1931 = opB[19] & opA[31];
logic p2000;
assign p2000 = opB[20] & opA[0];
logic p2001;
assign p2001 = opB[20] & opA[1];
logic p2002;
assign p2002 = opB[20] & opA[2];
logic p2003;
assign p2003 = opB[20] & opA[3];
logic p2004;
assign p2004 = opB[20] & opA[4];
logic p2005;
assign p2005 = opB[20] & opA[5];
logic p2006;
assign p2006 = opB[20] & opA[6];
logic p2007;
assign p2007 = opB[20] & opA[7];
logic p2008;
assign p2008 = opB[20] & opA[8];
logic p2009;
assign p2009 = opB[20] & opA[9];
logic p2010;
assign p2010 = opB[20] & opA[10];
logic p2011;
assign p2011 = opB[20] & opA[11];
logic p2012;
assign p2012 = opB[20] & opA[12];
logic p2013;
assign p2013 = opB[20] & opA[13];
logic p2014;
assign p2014 = opB[20] & opA[14];
logic p2015;
assign p2015 = opB[20] & opA[15];
logic p2016;
assign p2016 = opB[20] & opA[16];
logic p2017;
assign p2017 = opB[20] & opA[17];
logic p2018;
assign p2018 = opB[20] & opA[18];
logic p2019;
assign p2019 = opB[20] & opA[19];
logic p2020;
assign p2020 = opB[20] & opA[20];
logic p2021;
assign p2021 = opB[20] & opA[21];
logic p2022;
assign p2022 = opB[20] & opA[22];
logic p2023;
assign p2023 = opB[20] & opA[23];
logic p2024;
assign p2024 = opB[20] & opA[24];
logic p2025;
assign p2025 = opB[20] & opA[25];
logic p2026;
assign p2026 = opB[20] & opA[26];
logic p2027;
assign p2027 = opB[20] & opA[27];
logic p2028;
assign p2028 = opB[20] & opA[28];
logic p2029;
assign p2029 = opB[20] & opA[29];
logic p2030;
assign p2030 = opB[20] & opA[30];
logic p2031;
assign p2031 = opB[20] & opA[31];
logic p2100;
assign p2100 = opB[21] & opA[0];
logic p2101;
assign p2101 = opB[21] & opA[1];
logic p2102;
assign p2102 = opB[21] & opA[2];
logic p2103;
assign p2103 = opB[21] & opA[3];
logic p2104;
assign p2104 = opB[21] & opA[4];
logic p2105;
assign p2105 = opB[21] & opA[5];
logic p2106;
assign p2106 = opB[21] & opA[6];
logic p2107;
assign p2107 = opB[21] & opA[7];
logic p2108;
assign p2108 = opB[21] & opA[8];
logic p2109;
assign p2109 = opB[21] & opA[9];
logic p2110;
assign p2110 = opB[21] & opA[10];
logic p2111;
assign p2111 = opB[21] & opA[11];
logic p2112;
assign p2112 = opB[21] & opA[12];
logic p2113;
assign p2113 = opB[21] & opA[13];
logic p2114;
assign p2114 = opB[21] & opA[14];
logic p2115;
assign p2115 = opB[21] & opA[15];
logic p2116;
assign p2116 = opB[21] & opA[16];
logic p2117;
assign p2117 = opB[21] & opA[17];
logic p2118;
assign p2118 = opB[21] & opA[18];
logic p2119;
assign p2119 = opB[21] & opA[19];
logic p2120;
assign p2120 = opB[21] & opA[20];
logic p2121;
assign p2121 = opB[21] & opA[21];
logic p2122;
assign p2122 = opB[21] & opA[22];
logic p2123;
assign p2123 = opB[21] & opA[23];
logic p2124;
assign p2124 = opB[21] & opA[24];
logic p2125;
assign p2125 = opB[21] & opA[25];
logic p2126;
assign p2126 = opB[21] & opA[26];
logic p2127;
assign p2127 = opB[21] & opA[27];
logic p2128;
assign p2128 = opB[21] & opA[28];
logic p2129;
assign p2129 = opB[21] & opA[29];
logic p2130;
assign p2130 = opB[21] & opA[30];
logic p2131;
assign p2131 = opB[21] & opA[31];
logic p2200;
assign p2200 = opB[22] & opA[0];
logic p2201;
assign p2201 = opB[22] & opA[1];
logic p2202;
assign p2202 = opB[22] & opA[2];
logic p2203;
assign p2203 = opB[22] & opA[3];
logic p2204;
assign p2204 = opB[22] & opA[4];
logic p2205;
assign p2205 = opB[22] & opA[5];
logic p2206;
assign p2206 = opB[22] & opA[6];
logic p2207;
assign p2207 = opB[22] & opA[7];
logic p2208;
assign p2208 = opB[22] & opA[8];
logic p2209;
assign p2209 = opB[22] & opA[9];
logic p2210;
assign p2210 = opB[22] & opA[10];
logic p2211;
assign p2211 = opB[22] & opA[11];
logic p2212;
assign p2212 = opB[22] & opA[12];
logic p2213;
assign p2213 = opB[22] & opA[13];
logic p2214;
assign p2214 = opB[22] & opA[14];
logic p2215;
assign p2215 = opB[22] & opA[15];
logic p2216;
assign p2216 = opB[22] & opA[16];
logic p2217;
assign p2217 = opB[22] & opA[17];
logic p2218;
assign p2218 = opB[22] & opA[18];
logic p2219;
assign p2219 = opB[22] & opA[19];
logic p2220;
assign p2220 = opB[22] & opA[20];
logic p2221;
assign p2221 = opB[22] & opA[21];
logic p2222;
assign p2222 = opB[22] & opA[22];
logic p2223;
assign p2223 = opB[22] & opA[23];
logic p2224;
assign p2224 = opB[22] & opA[24];
logic p2225;
assign p2225 = opB[22] & opA[25];
logic p2226;
assign p2226 = opB[22] & opA[26];
logic p2227;
assign p2227 = opB[22] & opA[27];
logic p2228;
assign p2228 = opB[22] & opA[28];
logic p2229;
assign p2229 = opB[22] & opA[29];
logic p2230;
assign p2230 = opB[22] & opA[30];
logic p2231;
assign p2231 = opB[22] & opA[31];
logic p2300;
assign p2300 = opB[23] & opA[0];
logic p2301;
assign p2301 = opB[23] & opA[1];
logic p2302;
assign p2302 = opB[23] & opA[2];
logic p2303;
assign p2303 = opB[23] & opA[3];
logic p2304;
assign p2304 = opB[23] & opA[4];
logic p2305;
assign p2305 = opB[23] & opA[5];
logic p2306;
assign p2306 = opB[23] & opA[6];
logic p2307;
assign p2307 = opB[23] & opA[7];
logic p2308;
assign p2308 = opB[23] & opA[8];
logic p2309;
assign p2309 = opB[23] & opA[9];
logic p2310;
assign p2310 = opB[23] & opA[10];
logic p2311;
assign p2311 = opB[23] & opA[11];
logic p2312;
assign p2312 = opB[23] & opA[12];
logic p2313;
assign p2313 = opB[23] & opA[13];
logic p2314;
assign p2314 = opB[23] & opA[14];
logic p2315;
assign p2315 = opB[23] & opA[15];
logic p2316;
assign p2316 = opB[23] & opA[16];
logic p2317;
assign p2317 = opB[23] & opA[17];
logic p2318;
assign p2318 = opB[23] & opA[18];
logic p2319;
assign p2319 = opB[23] & opA[19];
logic p2320;
assign p2320 = opB[23] & opA[20];
logic p2321;
assign p2321 = opB[23] & opA[21];
logic p2322;
assign p2322 = opB[23] & opA[22];
logic p2323;
assign p2323 = opB[23] & opA[23];
logic p2324;
assign p2324 = opB[23] & opA[24];
logic p2325;
assign p2325 = opB[23] & opA[25];
logic p2326;
assign p2326 = opB[23] & opA[26];
logic p2327;
assign p2327 = opB[23] & opA[27];
logic p2328;
assign p2328 = opB[23] & opA[28];
logic p2329;
assign p2329 = opB[23] & opA[29];
logic p2330;
assign p2330 = opB[23] & opA[30];
logic p2331;
assign p2331 = opB[23] & opA[31];
logic p2400;
assign p2400 = opB[24] & opA[0];
logic p2401;
assign p2401 = opB[24] & opA[1];
logic p2402;
assign p2402 = opB[24] & opA[2];
logic p2403;
assign p2403 = opB[24] & opA[3];
logic p2404;
assign p2404 = opB[24] & opA[4];
logic p2405;
assign p2405 = opB[24] & opA[5];
logic p2406;
assign p2406 = opB[24] & opA[6];
logic p2407;
assign p2407 = opB[24] & opA[7];
logic p2408;
assign p2408 = opB[24] & opA[8];
logic p2409;
assign p2409 = opB[24] & opA[9];
logic p2410;
assign p2410 = opB[24] & opA[10];
logic p2411;
assign p2411 = opB[24] & opA[11];
logic p2412;
assign p2412 = opB[24] & opA[12];
logic p2413;
assign p2413 = opB[24] & opA[13];
logic p2414;
assign p2414 = opB[24] & opA[14];
logic p2415;
assign p2415 = opB[24] & opA[15];
logic p2416;
assign p2416 = opB[24] & opA[16];
logic p2417;
assign p2417 = opB[24] & opA[17];
logic p2418;
assign p2418 = opB[24] & opA[18];
logic p2419;
assign p2419 = opB[24] & opA[19];
logic p2420;
assign p2420 = opB[24] & opA[20];
logic p2421;
assign p2421 = opB[24] & opA[21];
logic p2422;
assign p2422 = opB[24] & opA[22];
logic p2423;
assign p2423 = opB[24] & opA[23];
logic p2424;
assign p2424 = opB[24] & opA[24];
logic p2425;
assign p2425 = opB[24] & opA[25];
logic p2426;
assign p2426 = opB[24] & opA[26];
logic p2427;
assign p2427 = opB[24] & opA[27];
logic p2428;
assign p2428 = opB[24] & opA[28];
logic p2429;
assign p2429 = opB[24] & opA[29];
logic p2430;
assign p2430 = opB[24] & opA[30];
logic p2431;
assign p2431 = opB[24] & opA[31];
logic p2500;
assign p2500 = opB[25] & opA[0];
logic p2501;
assign p2501 = opB[25] & opA[1];
logic p2502;
assign p2502 = opB[25] & opA[2];
logic p2503;
assign p2503 = opB[25] & opA[3];
logic p2504;
assign p2504 = opB[25] & opA[4];
logic p2505;
assign p2505 = opB[25] & opA[5];
logic p2506;
assign p2506 = opB[25] & opA[6];
logic p2507;
assign p2507 = opB[25] & opA[7];
logic p2508;
assign p2508 = opB[25] & opA[8];
logic p2509;
assign p2509 = opB[25] & opA[9];
logic p2510;
assign p2510 = opB[25] & opA[10];
logic p2511;
assign p2511 = opB[25] & opA[11];
logic p2512;
assign p2512 = opB[25] & opA[12];
logic p2513;
assign p2513 = opB[25] & opA[13];
logic p2514;
assign p2514 = opB[25] & opA[14];
logic p2515;
assign p2515 = opB[25] & opA[15];
logic p2516;
assign p2516 = opB[25] & opA[16];
logic p2517;
assign p2517 = opB[25] & opA[17];
logic p2518;
assign p2518 = opB[25] & opA[18];
logic p2519;
assign p2519 = opB[25] & opA[19];
logic p2520;
assign p2520 = opB[25] & opA[20];
logic p2521;
assign p2521 = opB[25] & opA[21];
logic p2522;
assign p2522 = opB[25] & opA[22];
logic p2523;
assign p2523 = opB[25] & opA[23];
logic p2524;
assign p2524 = opB[25] & opA[24];
logic p2525;
assign p2525 = opB[25] & opA[25];
logic p2526;
assign p2526 = opB[25] & opA[26];
logic p2527;
assign p2527 = opB[25] & opA[27];
logic p2528;
assign p2528 = opB[25] & opA[28];
logic p2529;
assign p2529 = opB[25] & opA[29];
logic p2530;
assign p2530 = opB[25] & opA[30];
logic p2531;
assign p2531 = opB[25] & opA[31];
logic p2600;
assign p2600 = opB[26] & opA[0];
logic p2601;
assign p2601 = opB[26] & opA[1];
logic p2602;
assign p2602 = opB[26] & opA[2];
logic p2603;
assign p2603 = opB[26] & opA[3];
logic p2604;
assign p2604 = opB[26] & opA[4];
logic p2605;
assign p2605 = opB[26] & opA[5];
logic p2606;
assign p2606 = opB[26] & opA[6];
logic p2607;
assign p2607 = opB[26] & opA[7];
logic p2608;
assign p2608 = opB[26] & opA[8];
logic p2609;
assign p2609 = opB[26] & opA[9];
logic p2610;
assign p2610 = opB[26] & opA[10];
logic p2611;
assign p2611 = opB[26] & opA[11];
logic p2612;
assign p2612 = opB[26] & opA[12];
logic p2613;
assign p2613 = opB[26] & opA[13];
logic p2614;
assign p2614 = opB[26] & opA[14];
logic p2615;
assign p2615 = opB[26] & opA[15];
logic p2616;
assign p2616 = opB[26] & opA[16];
logic p2617;
assign p2617 = opB[26] & opA[17];
logic p2618;
assign p2618 = opB[26] & opA[18];
logic p2619;
assign p2619 = opB[26] & opA[19];
logic p2620;
assign p2620 = opB[26] & opA[20];
logic p2621;
assign p2621 = opB[26] & opA[21];
logic p2622;
assign p2622 = opB[26] & opA[22];
logic p2623;
assign p2623 = opB[26] & opA[23];
logic p2624;
assign p2624 = opB[26] & opA[24];
logic p2625;
assign p2625 = opB[26] & opA[25];
logic p2626;
assign p2626 = opB[26] & opA[26];
logic p2627;
assign p2627 = opB[26] & opA[27];
logic p2628;
assign p2628 = opB[26] & opA[28];
logic p2629;
assign p2629 = opB[26] & opA[29];
logic p2630;
assign p2630 = opB[26] & opA[30];
logic p2631;
assign p2631 = opB[26] & opA[31];
logic p2700;
assign p2700 = opB[27] & opA[0];
logic p2701;
assign p2701 = opB[27] & opA[1];
logic p2702;
assign p2702 = opB[27] & opA[2];
logic p2703;
assign p2703 = opB[27] & opA[3];
logic p2704;
assign p2704 = opB[27] & opA[4];
logic p2705;
assign p2705 = opB[27] & opA[5];
logic p2706;
assign p2706 = opB[27] & opA[6];
logic p2707;
assign p2707 = opB[27] & opA[7];
logic p2708;
assign p2708 = opB[27] & opA[8];
logic p2709;
assign p2709 = opB[27] & opA[9];
logic p2710;
assign p2710 = opB[27] & opA[10];
logic p2711;
assign p2711 = opB[27] & opA[11];
logic p2712;
assign p2712 = opB[27] & opA[12];
logic p2713;
assign p2713 = opB[27] & opA[13];
logic p2714;
assign p2714 = opB[27] & opA[14];
logic p2715;
assign p2715 = opB[27] & opA[15];
logic p2716;
assign p2716 = opB[27] & opA[16];
logic p2717;
assign p2717 = opB[27] & opA[17];
logic p2718;
assign p2718 = opB[27] & opA[18];
logic p2719;
assign p2719 = opB[27] & opA[19];
logic p2720;
assign p2720 = opB[27] & opA[20];
logic p2721;
assign p2721 = opB[27] & opA[21];
logic p2722;
assign p2722 = opB[27] & opA[22];
logic p2723;
assign p2723 = opB[27] & opA[23];
logic p2724;
assign p2724 = opB[27] & opA[24];
logic p2725;
assign p2725 = opB[27] & opA[25];
logic p2726;
assign p2726 = opB[27] & opA[26];
logic p2727;
assign p2727 = opB[27] & opA[27];
logic p2728;
assign p2728 = opB[27] & opA[28];
logic p2729;
assign p2729 = opB[27] & opA[29];
logic p2730;
assign p2730 = opB[27] & opA[30];
logic p2731;
assign p2731 = opB[27] & opA[31];
logic p2800;
assign p2800 = opB[28] & opA[0];
logic p2801;
assign p2801 = opB[28] & opA[1];
logic p2802;
assign p2802 = opB[28] & opA[2];
logic p2803;
assign p2803 = opB[28] & opA[3];
logic p2804;
assign p2804 = opB[28] & opA[4];
logic p2805;
assign p2805 = opB[28] & opA[5];
logic p2806;
assign p2806 = opB[28] & opA[6];
logic p2807;
assign p2807 = opB[28] & opA[7];
logic p2808;
assign p2808 = opB[28] & opA[8];
logic p2809;
assign p2809 = opB[28] & opA[9];
logic p2810;
assign p2810 = opB[28] & opA[10];
logic p2811;
assign p2811 = opB[28] & opA[11];
logic p2812;
assign p2812 = opB[28] & opA[12];
logic p2813;
assign p2813 = opB[28] & opA[13];
logic p2814;
assign p2814 = opB[28] & opA[14];
logic p2815;
assign p2815 = opB[28] & opA[15];
logic p2816;
assign p2816 = opB[28] & opA[16];
logic p2817;
assign p2817 = opB[28] & opA[17];
logic p2818;
assign p2818 = opB[28] & opA[18];
logic p2819;
assign p2819 = opB[28] & opA[19];
logic p2820;
assign p2820 = opB[28] & opA[20];
logic p2821;
assign p2821 = opB[28] & opA[21];
logic p2822;
assign p2822 = opB[28] & opA[22];
logic p2823;
assign p2823 = opB[28] & opA[23];
logic p2824;
assign p2824 = opB[28] & opA[24];
logic p2825;
assign p2825 = opB[28] & opA[25];
logic p2826;
assign p2826 = opB[28] & opA[26];
logic p2827;
assign p2827 = opB[28] & opA[27];
logic p2828;
assign p2828 = opB[28] & opA[28];
logic p2829;
assign p2829 = opB[28] & opA[29];
logic p2830;
assign p2830 = opB[28] & opA[30];
logic p2831;
assign p2831 = opB[28] & opA[31];
logic p2900;
assign p2900 = opB[29] & opA[0];
logic p2901;
assign p2901 = opB[29] & opA[1];
logic p2902;
assign p2902 = opB[29] & opA[2];
logic p2903;
assign p2903 = opB[29] & opA[3];
logic p2904;
assign p2904 = opB[29] & opA[4];
logic p2905;
assign p2905 = opB[29] & opA[5];
logic p2906;
assign p2906 = opB[29] & opA[6];
logic p2907;
assign p2907 = opB[29] & opA[7];
logic p2908;
assign p2908 = opB[29] & opA[8];
logic p2909;
assign p2909 = opB[29] & opA[9];
logic p2910;
assign p2910 = opB[29] & opA[10];
logic p2911;
assign p2911 = opB[29] & opA[11];
logic p2912;
assign p2912 = opB[29] & opA[12];
logic p2913;
assign p2913 = opB[29] & opA[13];
logic p2914;
assign p2914 = opB[29] & opA[14];
logic p2915;
assign p2915 = opB[29] & opA[15];
logic p2916;
assign p2916 = opB[29] & opA[16];
logic p2917;
assign p2917 = opB[29] & opA[17];
logic p2918;
assign p2918 = opB[29] & opA[18];
logic p2919;
assign p2919 = opB[29] & opA[19];
logic p2920;
assign p2920 = opB[29] & opA[20];
logic p2921;
assign p2921 = opB[29] & opA[21];
logic p2922;
assign p2922 = opB[29] & opA[22];
logic p2923;
assign p2923 = opB[29] & opA[23];
logic p2924;
assign p2924 = opB[29] & opA[24];
logic p2925;
assign p2925 = opB[29] & opA[25];
logic p2926;
assign p2926 = opB[29] & opA[26];
logic p2927;
assign p2927 = opB[29] & opA[27];
logic p2928;
assign p2928 = opB[29] & opA[28];
logic p2929;
assign p2929 = opB[29] & opA[29];
logic p2930;
assign p2930 = opB[29] & opA[30];
logic p2931;
assign p2931 = opB[29] & opA[31];
logic p3000;
assign p3000 = opB[30] & opA[0];
logic p3001;
assign p3001 = opB[30] & opA[1];
logic p3002;
assign p3002 = opB[30] & opA[2];
logic p3003;
assign p3003 = opB[30] & opA[3];
logic p3004;
assign p3004 = opB[30] & opA[4];
logic p3005;
assign p3005 = opB[30] & opA[5];
logic p3006;
assign p3006 = opB[30] & opA[6];
logic p3007;
assign p3007 = opB[30] & opA[7];
logic p3008;
assign p3008 = opB[30] & opA[8];
logic p3009;
assign p3009 = opB[30] & opA[9];
logic p3010;
assign p3010 = opB[30] & opA[10];
logic p3011;
assign p3011 = opB[30] & opA[11];
logic p3012;
assign p3012 = opB[30] & opA[12];
logic p3013;
assign p3013 = opB[30] & opA[13];
logic p3014;
assign p3014 = opB[30] & opA[14];
logic p3015;
assign p3015 = opB[30] & opA[15];
logic p3016;
assign p3016 = opB[30] & opA[16];
logic p3017;
assign p3017 = opB[30] & opA[17];
logic p3018;
assign p3018 = opB[30] & opA[18];
logic p3019;
assign p3019 = opB[30] & opA[19];
logic p3020;
assign p3020 = opB[30] & opA[20];
logic p3021;
assign p3021 = opB[30] & opA[21];
logic p3022;
assign p3022 = opB[30] & opA[22];
logic p3023;
assign p3023 = opB[30] & opA[23];
logic p3024;
assign p3024 = opB[30] & opA[24];
logic p3025;
assign p3025 = opB[30] & opA[25];
logic p3026;
assign p3026 = opB[30] & opA[26];
logic p3027;
assign p3027 = opB[30] & opA[27];
logic p3028;
assign p3028 = opB[30] & opA[28];
logic p3029;
assign p3029 = opB[30] & opA[29];
logic p3030;
assign p3030 = opB[30] & opA[30];
logic p3031;
assign p3031 = opB[30] & opA[31];
logic p3100;
assign p3100 = opB[31] & opA[0];
logic p3101;
assign p3101 = opB[31] & opA[1];
logic p3102;
assign p3102 = opB[31] & opA[2];
logic p3103;
assign p3103 = opB[31] & opA[3];
logic p3104;
assign p3104 = opB[31] & opA[4];
logic p3105;
assign p3105 = opB[31] & opA[5];
logic p3106;
assign p3106 = opB[31] & opA[6];
logic p3107;
assign p3107 = opB[31] & opA[7];
logic p3108;
assign p3108 = opB[31] & opA[8];
logic p3109;
assign p3109 = opB[31] & opA[9];
logic p3110;
assign p3110 = opB[31] & opA[10];
logic p3111;
assign p3111 = opB[31] & opA[11];
logic p3112;
assign p3112 = opB[31] & opA[12];
logic p3113;
assign p3113 = opB[31] & opA[13];
logic p3114;
assign p3114 = opB[31] & opA[14];
logic p3115;
assign p3115 = opB[31] & opA[15];
logic p3116;
assign p3116 = opB[31] & opA[16];
logic p3117;
assign p3117 = opB[31] & opA[17];
logic p3118;
assign p3118 = opB[31] & opA[18];
logic p3119;
assign p3119 = opB[31] & opA[19];
logic p3120;
assign p3120 = opB[31] & opA[20];
logic p3121;
assign p3121 = opB[31] & opA[21];
logic p3122;
assign p3122 = opB[31] & opA[22];
logic p3123;
assign p3123 = opB[31] & opA[23];
logic p3124;
assign p3124 = opB[31] & opA[24];
logic p3125;
assign p3125 = opB[31] & opA[25];
logic p3126;
assign p3126 = opB[31] & opA[26];
logic p3127;
assign p3127 = opB[31] & opA[27];
logic p3128;
assign p3128 = opB[31] & opA[28];
logic p3129;
assign p3129 = opB[31] & opA[29];
logic p3130;
assign p3130 = opB[31] & opA[30];
logic p3131;
assign p3131 = opB[31] & opA[31];
// stage 8 begin ======================================================================= 
HA HA_s8_280(.A(comb[0][28]), .B(comb[1][27]), .S(S_s8_280), .c_out(C_s8_280));
FA FA_s8_290(.A(comb[0][29]), .B(comb[1][28]), .c_in(comb[2][27]), .S(S_s8_290), .c_out(C_s8_290));
HA HA_s8_291(.A(comb[3][26]), .B(comb[4][25]), .S(S_s8_291), .c_out(C_s8_291));
FA FA_s8_300(.A(comb[0][30]), .B(comb[1][29]), .c_in(comb[2][28]), .S(S_s8_300), .c_out(C_s8_300));
FA FA_s8_301(.A(comb[3][27]), .B(comb[4][26]), .c_in(comb[5][25]), .S(S_s8_301), .c_out(C_s8_301));
HA HA_s8_302(.A(comb[6][24]), .B(comb[7][23]), .S(S_s8_302), .c_out(C_s8_302));
FA FA_s8_310(.A(comb[0][31]), .B(comb[1][30]), .c_in(comb[2][29]), .S(S_s8_310), .c_out(C_s8_310));
FA FA_s8_311(.A(comb[3][28]), .B(comb[4][27]), .c_in(comb[5][26]), .S(S_s8_311), .c_out(C_s8_311));
FA FA_s8_312(.A(comb[6][25]), .B(comb[7][24]), .c_in(comb[8][23]), .S(S_s8_312), .c_out(C_s8_312));
HA HA_s8_313(.A(comb[9][22]), .B(comb[10][21]), .S(S_s8_313), .c_out(C_s8_313));
FA FA_s8_320(.A(comb[1][31]), .B(comb[2][30]), .c_in(comb[3][29]), .S(S_s8_320), .c_out(C_s8_320));
FA FA_s8_321(.A(comb[4][28]), .B(comb[5][27]), .c_in(comb[6][26]), .S(S_s8_321), .c_out(C_s8_321));
FA FA_s8_322(.A(comb[7][25]), .B(comb[8][24]), .c_in(comb[9][23]), .S(S_s8_322), .c_out(C_s8_322));
HA HA_s8_323(.A(comb[10][22]), .B(comb[11][21]), .S(S_s8_323), .c_out(C_s8_323));
FA FA_s8_330(.A(comb[2][31]), .B(comb[3][30]), .c_in(comb[4][29]), .S(S_s8_330), .c_out(C_s8_330));
FA FA_s8_331(.A(comb[5][28]), .B(comb[6][27]), .c_in(comb[7][26]), .S(S_s8_331), .c_out(C_s8_331));
FA FA_s8_332(.A(comb[8][25]), .B(comb[9][24]), .c_in(comb[10][23]), .S(S_s8_332), .c_out(C_s8_332));
FA FA_s8_340(.A(comb[3][31]), .B(comb[4][30]), .c_in(comb[5][29]), .S(S_s8_340), .c_out(C_s8_340));
FA FA_s8_341(.A(comb[6][28]), .B(comb[7][27]), .c_in(comb[8][26]), .S(S_s8_341), .c_out(C_s8_341));
FA FA_s8_350(.A(comb[4][31]), .B(comb[5][30]), .c_in(comb[6][29]), .S(S_s8_350), .c_out(C_s8_350));
// stage 8 end ======================================================================= 

// stage 7 begin ======================================================================= 
HA HA_s7_190(.A(comb[0][19]), .B(comb[1][18]), .S(S_s7_190), .c_out(C_s7_190));
FA FA_s7_200(.A(comb[0][20]), .B(comb[1][19]), .c_in(comb[2][18]), .S(S_s7_200), .c_out(C_s7_200));
HA HA_s7_201(.A(comb[3][17]), .B(comb[4][16]), .S(S_s7_201), .c_out(C_s7_201));
FA FA_s7_210(.A(comb[0][21]), .B(comb[1][20]), .c_in(comb[2][19]), .S(S_s7_210), .c_out(C_s7_210));
FA FA_s7_211(.A(comb[3][18]), .B(comb[4][17]), .c_in(comb[5][16]), .S(S_s7_211), .c_out(C_s7_211));
HA HA_s7_212(.A(comb[6][15]), .B(comb[7][14]), .S(S_s7_212), .c_out(C_s7_212));
FA FA_s7_220(.A(comb[0][22]), .B(comb[1][21]), .c_in(comb[2][20]), .S(S_s7_220), .c_out(C_s7_220));
FA FA_s7_221(.A(comb[3][19]), .B(comb[4][18]), .c_in(comb[5][17]), .S(S_s7_221), .c_out(C_s7_221));
FA FA_s7_222(.A(comb[6][16]), .B(comb[7][15]), .c_in(comb[8][14]), .S(S_s7_222), .c_out(C_s7_222));
HA HA_s7_223(.A(comb[9][13]), .B(comb[10][12]), .S(S_s7_223), .c_out(C_s7_223));
FA FA_s7_230(.A(comb[0][23]), .B(comb[1][22]), .c_in(comb[2][21]), .S(S_s7_230), .c_out(C_s7_230));
FA FA_s7_231(.A(comb[3][20]), .B(comb[4][19]), .c_in(comb[5][18]), .S(S_s7_231), .c_out(C_s7_231));
FA FA_s7_232(.A(comb[6][17]), .B(comb[7][16]), .c_in(comb[8][15]), .S(S_s7_232), .c_out(C_s7_232));
FA FA_s7_233(.A(comb[9][14]), .B(comb[10][13]), .c_in(comb[11][12]), .S(S_s7_233), .c_out(C_s7_233));
HA HA_s7_234(.A(comb[12][11]), .B(comb[13][10]), .S(S_s7_234), .c_out(C_s7_234));
FA FA_s7_240(.A(comb[0][24]), .B(comb[1][23]), .c_in(comb[2][22]), .S(S_s7_240), .c_out(C_s7_240));
FA FA_s7_241(.A(comb[3][21]), .B(comb[4][20]), .c_in(comb[5][19]), .S(S_s7_241), .c_out(C_s7_241));
FA FA_s7_242(.A(comb[6][18]), .B(comb[7][17]), .c_in(comb[8][16]), .S(S_s7_242), .c_out(C_s7_242));
FA FA_s7_243(.A(comb[9][15]), .B(comb[10][14]), .c_in(comb[11][13]), .S(S_s7_243), .c_out(C_s7_243));
FA FA_s7_244(.A(comb[12][12]), .B(comb[13][11]), .c_in(comb[14][10]), .S(S_s7_244), .c_out(C_s7_244));
HA HA_s7_245(.A(comb[15][9]), .B(comb[16][8]), .S(S_s7_245), .c_out(C_s7_245));
FA FA_s7_250(.A(comb[0][25]), .B(comb[1][24]), .c_in(comb[2][23]), .S(S_s7_250), .c_out(C_s7_250));
FA FA_s7_251(.A(comb[3][22]), .B(comb[4][21]), .c_in(comb[5][20]), .S(S_s7_251), .c_out(C_s7_251));
FA FA_s7_252(.A(comb[6][19]), .B(comb[7][18]), .c_in(comb[8][17]), .S(S_s7_252), .c_out(C_s7_252));
FA FA_s7_253(.A(comb[9][16]), .B(comb[10][15]), .c_in(comb[11][14]), .S(S_s7_253), .c_out(C_s7_253));
FA FA_s7_254(.A(comb[12][13]), .B(comb[13][12]), .c_in(comb[14][11]), .S(S_s7_254), .c_out(C_s7_254));
FA FA_s7_255(.A(comb[15][10]), .B(comb[16][9]), .c_in(comb[17][8]), .S(S_s7_255), .c_out(C_s7_255));
HA HA_s7_256(.A(comb[18][7]), .B(comb[19][6]), .S(S_s7_256), .c_out(C_s7_256));
FA FA_s7_260(.A(comb[0][26]), .B(comb[1][25]), .c_in(comb[2][24]), .S(S_s7_260), .c_out(C_s7_260));
FA FA_s7_261(.A(comb[3][23]), .B(comb[4][22]), .c_in(comb[5][21]), .S(S_s7_261), .c_out(C_s7_261));
FA FA_s7_262(.A(comb[6][20]), .B(comb[7][19]), .c_in(comb[8][18]), .S(S_s7_262), .c_out(C_s7_262));
FA FA_s7_263(.A(comb[9][17]), .B(comb[10][16]), .c_in(comb[11][15]), .S(S_s7_263), .c_out(C_s7_263));
FA FA_s7_264(.A(comb[12][14]), .B(comb[13][13]), .c_in(comb[14][12]), .S(S_s7_264), .c_out(C_s7_264));
FA FA_s7_265(.A(comb[15][11]), .B(comb[16][10]), .c_in(comb[17][9]), .S(S_s7_265), .c_out(C_s7_265));
FA FA_s7_266(.A(comb[18][8]), .B(comb[19][7]), .c_in(comb[20][6]), .S(S_s7_266), .c_out(C_s7_266));
HA HA_s7_267(.A(comb[21][5]), .B(comb[22][4]), .S(S_s7_267), .c_out(C_s7_267));
FA FA_s7_270(.A(comb[0][27]), .B(comb[1][26]), .c_in(comb[2][25]), .S(S_s7_270), .c_out(C_s7_270));
FA FA_s7_271(.A(comb[3][24]), .B(comb[4][23]), .c_in(comb[5][22]), .S(S_s7_271), .c_out(C_s7_271));
FA FA_s7_272(.A(comb[6][21]), .B(comb[7][20]), .c_in(comb[8][19]), .S(S_s7_272), .c_out(C_s7_272));
FA FA_s7_273(.A(comb[9][18]), .B(comb[10][17]), .c_in(comb[11][16]), .S(S_s7_273), .c_out(C_s7_273));
FA FA_s7_274(.A(comb[12][15]), .B(comb[13][14]), .c_in(comb[14][13]), .S(S_s7_274), .c_out(C_s7_274));
FA FA_s7_275(.A(comb[15][12]), .B(comb[16][11]), .c_in(comb[17][10]), .S(S_s7_275), .c_out(C_s7_275));
FA FA_s7_276(.A(comb[18][9]), .B(comb[19][8]), .c_in(comb[20][7]), .S(S_s7_276), .c_out(C_s7_276));
FA FA_s7_277(.A(comb[21][6]), .B(comb[22][5]), .c_in(comb[23][4]), .S(S_s7_277), .c_out(C_s7_277));
HA HA_s7_278(.A(comb[24][3]), .B(comb[25][2]), .S(S_s7_278), .c_out(C_s7_278));
FA FA_s7_280(.A(S_s8_280), .B(comb[2][26]), .c_in(comb[3][25]), .S(S_s7_280), .c_out(C_s7_280));
FA FA_s7_281(.A(comb[4][24]), .B(comb[5][23]), .c_in(comb[6][22]), .S(S_s7_281), .c_out(C_s7_281));
FA FA_s7_282(.A(comb[7][21]), .B(comb[8][20]), .c_in(comb[9][19]), .S(S_s7_282), .c_out(C_s7_282));
FA FA_s7_283(.A(comb[10][18]), .B(comb[11][17]), .c_in(comb[12][16]), .S(S_s7_283), .c_out(C_s7_283));
FA FA_s7_284(.A(comb[13][15]), .B(comb[14][14]), .c_in(comb[15][13]), .S(S_s7_284), .c_out(C_s7_284));
FA FA_s7_285(.A(comb[16][12]), .B(comb[17][11]), .c_in(comb[18][10]), .S(S_s7_285), .c_out(C_s7_285));
FA FA_s7_286(.A(comb[19][9]), .B(comb[20][8]), .c_in(comb[21][7]), .S(S_s7_286), .c_out(C_s7_286));
FA FA_s7_287(.A(comb[22][6]), .B(comb[23][5]), .c_in(comb[24][4]), .S(S_s7_287), .c_out(C_s7_287));
FA FA_s7_288(.A(comb[25][3]), .B(comb[26][2]), .c_in(comb[27][1]), .S(S_s7_288), .c_out(C_s7_288));
FA FA_s7_290(.A(S_s8_291), .B(S_s8_290), .c_in(C_s8_280), .S(S_s7_290), .c_out(C_s7_290));
FA FA_s7_291(.A(comb[5][24]), .B(comb[6][23]), .c_in(comb[7][22]), .S(S_s7_291), .c_out(C_s7_291));
FA FA_s7_292(.A(comb[8][21]), .B(comb[9][20]), .c_in(comb[10][19]), .S(S_s7_292), .c_out(C_s7_292));
FA FA_s7_293(.A(comb[11][18]), .B(comb[12][17]), .c_in(comb[13][16]), .S(S_s7_293), .c_out(C_s7_293));
FA FA_s7_294(.A(comb[14][15]), .B(comb[15][14]), .c_in(comb[16][13]), .S(S_s7_294), .c_out(C_s7_294));
FA FA_s7_295(.A(comb[17][12]), .B(comb[18][11]), .c_in(comb[19][10]), .S(S_s7_295), .c_out(C_s7_295));
FA FA_s7_296(.A(comb[20][9]), .B(comb[21][8]), .c_in(comb[22][7]), .S(S_s7_296), .c_out(C_s7_296));
FA FA_s7_297(.A(comb[23][6]), .B(comb[24][5]), .c_in(comb[25][4]), .S(S_s7_297), .c_out(C_s7_297));
FA FA_s7_298(.A(comb[26][3]), .B(comb[27][2]), .c_in(comb[28][1]), .S(S_s7_298), .c_out(C_s7_298));
FA FA_s7_300(.A(S_s8_302), .B(S_s8_301), .c_in(S_s8_300), .S(S_s7_300), .c_out(C_s7_300));
FA FA_s7_301(.A(C_s8_291), .B(C_s8_290), .c_in(comb[8][22]), .S(S_s7_301), .c_out(C_s7_301));
FA FA_s7_302(.A(comb[9][21]), .B(comb[10][20]), .c_in(comb[11][19]), .S(S_s7_302), .c_out(C_s7_302));
FA FA_s7_303(.A(comb[12][18]), .B(comb[13][17]), .c_in(comb[14][16]), .S(S_s7_303), .c_out(C_s7_303));
FA FA_s7_304(.A(comb[15][15]), .B(comb[16][14]), .c_in(comb[17][13]), .S(S_s7_304), .c_out(C_s7_304));
FA FA_s7_305(.A(comb[18][12]), .B(comb[19][11]), .c_in(comb[20][10]), .S(S_s7_305), .c_out(C_s7_305));
FA FA_s7_306(.A(comb[21][9]), .B(comb[22][8]), .c_in(comb[23][7]), .S(S_s7_306), .c_out(C_s7_306));
FA FA_s7_307(.A(comb[24][6]), .B(comb[25][5]), .c_in(comb[26][4]), .S(S_s7_307), .c_out(C_s7_307));
FA FA_s7_308(.A(comb[27][3]), .B(comb[28][2]), .c_in(comb[29][1]), .S(S_s7_308), .c_out(C_s7_308));
FA FA_s7_310(.A(S_s8_313), .B(S_s8_312), .c_in(S_s8_311), .S(S_s7_310), .c_out(C_s7_310));
FA FA_s7_311(.A(S_s8_310), .B(C_s8_302), .c_in(C_s8_301), .S(S_s7_311), .c_out(C_s7_311));
FA FA_s7_312(.A(C_s8_300), .B(comb[11][20]), .c_in(comb[12][19]), .S(S_s7_312), .c_out(C_s7_312));
FA FA_s7_313(.A(comb[13][18]), .B(comb[14][17]), .c_in(comb[15][16]), .S(S_s7_313), .c_out(C_s7_313));
FA FA_s7_314(.A(comb[16][15]), .B(comb[17][14]), .c_in(comb[18][13]), .S(S_s7_314), .c_out(C_s7_314));
FA FA_s7_315(.A(comb[19][12]), .B(comb[20][11]), .c_in(comb[21][10]), .S(S_s7_315), .c_out(C_s7_315));
FA FA_s7_316(.A(comb[22][9]), .B(comb[23][8]), .c_in(comb[24][7]), .S(S_s7_316), .c_out(C_s7_316));
FA FA_s7_317(.A(comb[25][6]), .B(comb[26][5]), .c_in(comb[27][4]), .S(S_s7_317), .c_out(C_s7_317));
FA FA_s7_318(.A(comb[28][3]), .B(comb[29][2]), .c_in(comb[30][1]), .S(S_s7_318), .c_out(C_s7_318));
FA FA_s7_320(.A(S_s8_323), .B(S_s8_322), .c_in(S_s8_321), .S(S_s7_320), .c_out(C_s7_320));
FA FA_s7_321(.A(S_s8_320), .B(C_s8_313), .c_in(C_s8_312), .S(S_s7_321), .c_out(C_s7_321));
FA FA_s7_322(.A(C_s8_311), .B(C_s8_310), .c_in(comb[12][20]), .S(S_s7_322), .c_out(C_s7_322));
FA FA_s7_323(.A(comb[13][19]), .B(comb[14][18]), .c_in(comb[15][17]), .S(S_s7_323), .c_out(C_s7_323));
FA FA_s7_324(.A(comb[16][16]), .B(comb[17][15]), .c_in(comb[18][14]), .S(S_s7_324), .c_out(C_s7_324));
FA FA_s7_325(.A(comb[19][13]), .B(comb[20][12]), .c_in(comb[21][11]), .S(S_s7_325), .c_out(C_s7_325));
FA FA_s7_326(.A(comb[22][10]), .B(comb[23][9]), .c_in(comb[24][8]), .S(S_s7_326), .c_out(C_s7_326));
FA FA_s7_327(.A(comb[25][7]), .B(comb[26][6]), .c_in(comb[27][5]), .S(S_s7_327), .c_out(C_s7_327));
FA FA_s7_328(.A(comb[28][4]), .B(comb[29][3]), .c_in(comb[30][2]), .S(S_s7_328), .c_out(C_s7_328));
FA FA_s7_330(.A(S_s8_332), .B(S_s8_331), .c_in(S_s8_330), .S(S_s7_330), .c_out(C_s7_330));
FA FA_s7_331(.A(C_s8_323), .B(C_s8_322), .c_in(C_s8_321), .S(S_s7_331), .c_out(C_s7_331));
FA FA_s7_332(.A(C_s8_320), .B(comb[11][22]), .c_in(comb[12][21]), .S(S_s7_332), .c_out(C_s7_332));
FA FA_s7_333(.A(comb[13][20]), .B(comb[14][19]), .c_in(comb[15][18]), .S(S_s7_333), .c_out(C_s7_333));
FA FA_s7_334(.A(comb[16][17]), .B(comb[17][16]), .c_in(comb[18][15]), .S(S_s7_334), .c_out(C_s7_334));
FA FA_s7_335(.A(comb[19][14]), .B(comb[20][13]), .c_in(comb[21][12]), .S(S_s7_335), .c_out(C_s7_335));
FA FA_s7_336(.A(comb[22][11]), .B(comb[23][10]), .c_in(comb[24][9]), .S(S_s7_336), .c_out(C_s7_336));
FA FA_s7_337(.A(comb[25][8]), .B(comb[26][7]), .c_in(comb[27][6]), .S(S_s7_337), .c_out(C_s7_337));
FA FA_s7_338(.A(comb[28][5]), .B(comb[29][4]), .c_in(comb[30][3]), .S(S_s7_338), .c_out(C_s7_338));
FA FA_s7_340(.A(S_s8_341), .B(S_s8_340), .c_in(C_s8_332), .S(S_s7_340), .c_out(C_s7_340));
FA FA_s7_341(.A(C_s8_331), .B(C_s8_330), .c_in(comb[9][25]), .S(S_s7_341), .c_out(C_s7_341));
FA FA_s7_342(.A(comb[10][24]), .B(comb[11][23]), .c_in(comb[12][22]), .S(S_s7_342), .c_out(C_s7_342));
FA FA_s7_343(.A(comb[13][21]), .B(comb[14][20]), .c_in(comb[15][19]), .S(S_s7_343), .c_out(C_s7_343));
FA FA_s7_344(.A(comb[16][18]), .B(comb[17][17]), .c_in(comb[18][16]), .S(S_s7_344), .c_out(C_s7_344));
FA FA_s7_345(.A(comb[19][15]), .B(comb[20][14]), .c_in(comb[21][13]), .S(S_s7_345), .c_out(C_s7_345));
FA FA_s7_346(.A(comb[22][12]), .B(comb[23][11]), .c_in(comb[24][10]), .S(S_s7_346), .c_out(C_s7_346));
FA FA_s7_347(.A(comb[25][9]), .B(comb[26][8]), .c_in(comb[27][7]), .S(S_s7_347), .c_out(C_s7_347));
FA FA_s7_348(.A(comb[28][6]), .B(comb[29][5]), .c_in(comb[30][4]), .S(S_s7_348), .c_out(C_s7_348));
FA FA_s7_350(.A(S_s8_350), .B(C_s8_341), .c_in(C_s8_340), .S(S_s7_350), .c_out(C_s7_350));
FA FA_s7_351(.A(comb[7][28]), .B(comb[8][27]), .c_in(comb[9][26]), .S(S_s7_351), .c_out(C_s7_351));
FA FA_s7_352(.A(comb[10][25]), .B(comb[11][24]), .c_in(comb[12][23]), .S(S_s7_352), .c_out(C_s7_352));
FA FA_s7_353(.A(comb[13][22]), .B(comb[14][21]), .c_in(comb[15][20]), .S(S_s7_353), .c_out(C_s7_353));
FA FA_s7_354(.A(comb[16][19]), .B(comb[17][18]), .c_in(comb[18][17]), .S(S_s7_354), .c_out(C_s7_354));
FA FA_s7_355(.A(comb[19][16]), .B(comb[20][15]), .c_in(comb[21][14]), .S(S_s7_355), .c_out(C_s7_355));
FA FA_s7_356(.A(comb[22][13]), .B(comb[23][12]), .c_in(comb[24][11]), .S(S_s7_356), .c_out(C_s7_356));
FA FA_s7_357(.A(comb[25][10]), .B(comb[26][9]), .c_in(comb[27][8]), .S(S_s7_357), .c_out(C_s7_357));
FA FA_s7_358(.A(comb[28][7]), .B(comb[29][6]), .c_in(comb[30][5]), .S(S_s7_358), .c_out(C_s7_358));
FA FA_s7_360(.A(C_s8_350), .B(comb[5][31]), .c_in(comb[6][30]), .S(S_s7_360), .c_out(C_s7_360));
FA FA_s7_361(.A(comb[7][29]), .B(comb[8][28]), .c_in(comb[9][27]), .S(S_s7_361), .c_out(C_s7_361));
FA FA_s7_362(.A(comb[10][26]), .B(comb[11][25]), .c_in(comb[12][24]), .S(S_s7_362), .c_out(C_s7_362));
FA FA_s7_363(.A(comb[13][23]), .B(comb[14][22]), .c_in(comb[15][21]), .S(S_s7_363), .c_out(C_s7_363));
FA FA_s7_364(.A(comb[16][20]), .B(comb[17][19]), .c_in(comb[18][18]), .S(S_s7_364), .c_out(C_s7_364));
FA FA_s7_365(.A(comb[19][17]), .B(comb[20][16]), .c_in(comb[21][15]), .S(S_s7_365), .c_out(C_s7_365));
FA FA_s7_366(.A(comb[22][14]), .B(comb[23][13]), .c_in(comb[24][12]), .S(S_s7_366), .c_out(C_s7_366));
FA FA_s7_367(.A(comb[25][11]), .B(comb[26][10]), .c_in(comb[27][9]), .S(S_s7_367), .c_out(C_s7_367));
FA FA_s7_368(.A(comb[28][8]), .B(comb[29][7]), .c_in(comb[30][6]), .S(S_s7_368), .c_out(C_s7_368));
FA FA_s7_370(.A(comb[6][31]), .B(comb[7][30]), .c_in(comb[8][29]), .S(S_s7_370), .c_out(C_s7_370));
FA FA_s7_371(.A(comb[9][28]), .B(comb[10][27]), .c_in(comb[11][26]), .S(S_s7_371), .c_out(C_s7_371));
FA FA_s7_372(.A(comb[12][25]), .B(comb[13][24]), .c_in(comb[14][23]), .S(S_s7_372), .c_out(C_s7_372));
FA FA_s7_373(.A(comb[15][22]), .B(comb[16][21]), .c_in(comb[17][20]), .S(S_s7_373), .c_out(C_s7_373));
FA FA_s7_374(.A(comb[18][19]), .B(comb[19][18]), .c_in(comb[20][17]), .S(S_s7_374), .c_out(C_s7_374));
FA FA_s7_375(.A(comb[21][16]), .B(comb[22][15]), .c_in(comb[23][14]), .S(S_s7_375), .c_out(C_s7_375));
FA FA_s7_376(.A(comb[24][13]), .B(comb[25][12]), .c_in(comb[26][11]), .S(S_s7_376), .c_out(C_s7_376));
FA FA_s7_377(.A(comb[27][10]), .B(comb[28][9]), .c_in(comb[29][8]), .S(S_s7_377), .c_out(C_s7_377));
FA FA_s7_380(.A(comb[7][31]), .B(comb[8][30]), .c_in(comb[9][29]), .S(S_s7_380), .c_out(C_s7_380));
FA FA_s7_381(.A(comb[10][28]), .B(comb[11][27]), .c_in(comb[12][26]), .S(S_s7_381), .c_out(C_s7_381));
FA FA_s7_382(.A(comb[13][25]), .B(comb[14][24]), .c_in(comb[15][23]), .S(S_s7_382), .c_out(C_s7_382));
FA FA_s7_383(.A(comb[16][22]), .B(comb[17][21]), .c_in(comb[18][20]), .S(S_s7_383), .c_out(C_s7_383));
FA FA_s7_384(.A(comb[19][19]), .B(comb[20][18]), .c_in(comb[21][17]), .S(S_s7_384), .c_out(C_s7_384));
FA FA_s7_385(.A(comb[22][16]), .B(comb[23][15]), .c_in(comb[24][14]), .S(S_s7_385), .c_out(C_s7_385));
FA FA_s7_386(.A(comb[25][13]), .B(comb[26][12]), .c_in(comb[27][11]), .S(S_s7_386), .c_out(C_s7_386));
FA FA_s7_390(.A(comb[8][31]), .B(comb[9][30]), .c_in(comb[10][29]), .S(S_s7_390), .c_out(C_s7_390));
FA FA_s7_391(.A(comb[11][28]), .B(comb[12][27]), .c_in(comb[13][26]), .S(S_s7_391), .c_out(C_s7_391));
FA FA_s7_392(.A(comb[14][25]), .B(comb[15][24]), .c_in(comb[16][23]), .S(S_s7_392), .c_out(C_s7_392));
FA FA_s7_393(.A(comb[17][22]), .B(comb[18][21]), .c_in(comb[19][20]), .S(S_s7_393), .c_out(C_s7_393));
FA FA_s7_394(.A(comb[20][19]), .B(comb[21][18]), .c_in(comb[22][17]), .S(S_s7_394), .c_out(C_s7_394));
FA FA_s7_395(.A(comb[23][16]), .B(comb[24][15]), .c_in(comb[25][14]), .S(S_s7_395), .c_out(C_s7_395));
FA FA_s7_400(.A(comb[9][31]), .B(comb[10][30]), .c_in(comb[11][29]), .S(S_s7_400), .c_out(C_s7_400));
FA FA_s7_401(.A(comb[12][28]), .B(comb[13][27]), .c_in(comb[14][26]), .S(S_s7_401), .c_out(C_s7_401));
FA FA_s7_402(.A(comb[15][25]), .B(comb[16][24]), .c_in(comb[17][23]), .S(S_s7_402), .c_out(C_s7_402));
FA FA_s7_403(.A(comb[18][22]), .B(comb[19][21]), .c_in(comb[20][20]), .S(S_s7_403), .c_out(C_s7_403));
FA FA_s7_404(.A(comb[21][19]), .B(comb[22][18]), .c_in(comb[23][17]), .S(S_s7_404), .c_out(C_s7_404));
FA FA_s7_410(.A(comb[10][31]), .B(comb[11][30]), .c_in(comb[12][29]), .S(S_s7_410), .c_out(C_s7_410));
FA FA_s7_411(.A(comb[13][28]), .B(comb[14][27]), .c_in(comb[15][26]), .S(S_s7_411), .c_out(C_s7_411));
FA FA_s7_412(.A(comb[16][25]), .B(comb[17][24]), .c_in(comb[18][23]), .S(S_s7_412), .c_out(C_s7_412));
FA FA_s7_413(.A(comb[19][22]), .B(comb[20][21]), .c_in(comb[21][20]), .S(S_s7_413), .c_out(C_s7_413));
FA FA_s7_420(.A(comb[11][31]), .B(comb[12][30]), .c_in(comb[13][29]), .S(S_s7_420), .c_out(C_s7_420));
FA FA_s7_421(.A(comb[14][28]), .B(comb[15][27]), .c_in(comb[16][26]), .S(S_s7_421), .c_out(C_s7_421));
FA FA_s7_422(.A(comb[17][25]), .B(comb[18][24]), .c_in(comb[19][23]), .S(S_s7_422), .c_out(C_s7_422));
FA FA_s7_430(.A(comb[12][31]), .B(comb[13][30]), .c_in(comb[14][29]), .S(S_s7_430), .c_out(C_s7_430));
FA FA_s7_431(.A(comb[15][28]), .B(comb[16][27]), .c_in(comb[17][26]), .S(S_s7_431), .c_out(C_s7_431));
FA FA_s7_440(.A(comb[13][31]), .B(comb[14][30]), .c_in(comb[15][29]), .S(S_s7_440), .c_out(C_s7_440));
// stage 7 end ======================================================================= 

// stage 6 begin ======================================================================= 
HA HA_s6_130(.A(comb[0][13]), .B(comb[1][12]), .S(S_s6_130), .c_out(C_s6_130));
FA FA_s6_140(.A(comb[0][14]), .B(comb[1][13]), .c_in(comb[2][12]), .S(S_s6_140), .c_out(C_s6_140));
HA HA_s6_141(.A(comb[3][11]), .B(comb[4][10]), .S(S_s6_141), .c_out(C_s6_141));
FA FA_s6_150(.A(comb[0][15]), .B(comb[1][14]), .c_in(comb[2][13]), .S(S_s6_150), .c_out(C_s6_150));
FA FA_s6_151(.A(comb[3][12]), .B(comb[4][11]), .c_in(comb[5][10]), .S(S_s6_151), .c_out(C_s6_151));
HA HA_s6_152(.A(comb[6][9]), .B(comb[7][8]), .S(S_s6_152), .c_out(C_s6_152));
FA FA_s6_160(.A(comb[0][16]), .B(comb[1][15]), .c_in(comb[2][14]), .S(S_s6_160), .c_out(C_s6_160));
FA FA_s6_161(.A(comb[3][13]), .B(comb[4][12]), .c_in(comb[5][11]), .S(S_s6_161), .c_out(C_s6_161));
FA FA_s6_162(.A(comb[6][10]), .B(comb[7][9]), .c_in(comb[8][8]), .S(S_s6_162), .c_out(C_s6_162));
HA HA_s6_163(.A(comb[9][7]), .B(comb[10][6]), .S(S_s6_163), .c_out(C_s6_163));
FA FA_s6_170(.A(comb[0][17]), .B(comb[1][16]), .c_in(comb[2][15]), .S(S_s6_170), .c_out(C_s6_170));
FA FA_s6_171(.A(comb[3][14]), .B(comb[4][13]), .c_in(comb[5][12]), .S(S_s6_171), .c_out(C_s6_171));
FA FA_s6_172(.A(comb[6][11]), .B(comb[7][10]), .c_in(comb[8][9]), .S(S_s6_172), .c_out(C_s6_172));
FA FA_s6_173(.A(comb[9][8]), .B(comb[10][7]), .c_in(comb[11][6]), .S(S_s6_173), .c_out(C_s6_173));
HA HA_s6_174(.A(comb[12][5]), .B(comb[13][4]), .S(S_s6_174), .c_out(C_s6_174));
FA FA_s6_180(.A(comb[0][18]), .B(comb[1][17]), .c_in(comb[2][16]), .S(S_s6_180), .c_out(C_s6_180));
FA FA_s6_181(.A(comb[3][15]), .B(comb[4][14]), .c_in(comb[5][13]), .S(S_s6_181), .c_out(C_s6_181));
FA FA_s6_182(.A(comb[6][12]), .B(comb[7][11]), .c_in(comb[8][10]), .S(S_s6_182), .c_out(C_s6_182));
FA FA_s6_183(.A(comb[9][9]), .B(comb[10][8]), .c_in(comb[11][7]), .S(S_s6_183), .c_out(C_s6_183));
FA FA_s6_184(.A(comb[12][6]), .B(comb[13][5]), .c_in(comb[14][4]), .S(S_s6_184), .c_out(C_s6_184));
HA HA_s6_185(.A(comb[15][3]), .B(comb[16][2]), .S(S_s6_185), .c_out(C_s6_185));
FA FA_s6_190(.A(S_s7_190), .B(comb[2][17]), .c_in(comb[3][16]), .S(S_s6_190), .c_out(C_s6_190));
FA FA_s6_191(.A(comb[4][15]), .B(comb[5][14]), .c_in(comb[6][13]), .S(S_s6_191), .c_out(C_s6_191));
FA FA_s6_192(.A(comb[7][12]), .B(comb[8][11]), .c_in(comb[9][10]), .S(S_s6_192), .c_out(C_s6_192));
FA FA_s6_193(.A(comb[10][9]), .B(comb[11][8]), .c_in(comb[12][7]), .S(S_s6_193), .c_out(C_s6_193));
FA FA_s6_194(.A(comb[13][6]), .B(comb[14][5]), .c_in(comb[15][4]), .S(S_s6_194), .c_out(C_s6_194));
FA FA_s6_195(.A(comb[16][3]), .B(comb[17][2]), .c_in(comb[18][1]), .S(S_s6_195), .c_out(C_s6_195));
FA FA_s6_200(.A(S_s7_201), .B(S_s7_200), .c_in(C_s7_190), .S(S_s6_200), .c_out(C_s6_200));
FA FA_s6_201(.A(comb[5][15]), .B(comb[6][14]), .c_in(comb[7][13]), .S(S_s6_201), .c_out(C_s6_201));
FA FA_s6_202(.A(comb[8][12]), .B(comb[9][11]), .c_in(comb[10][10]), .S(S_s6_202), .c_out(C_s6_202));
FA FA_s6_203(.A(comb[11][9]), .B(comb[12][8]), .c_in(comb[13][7]), .S(S_s6_203), .c_out(C_s6_203));
FA FA_s6_204(.A(comb[14][6]), .B(comb[15][5]), .c_in(comb[16][4]), .S(S_s6_204), .c_out(C_s6_204));
FA FA_s6_205(.A(comb[17][3]), .B(comb[18][2]), .c_in(comb[19][1]), .S(S_s6_205), .c_out(C_s6_205));
FA FA_s6_210(.A(S_s7_212), .B(S_s7_211), .c_in(S_s7_210), .S(S_s6_210), .c_out(C_s6_210));
FA FA_s6_211(.A(C_s7_201), .B(C_s7_200), .c_in(comb[8][13]), .S(S_s6_211), .c_out(C_s6_211));
FA FA_s6_212(.A(comb[9][12]), .B(comb[10][11]), .c_in(comb[11][10]), .S(S_s6_212), .c_out(C_s6_212));
FA FA_s6_213(.A(comb[12][9]), .B(comb[13][8]), .c_in(comb[14][7]), .S(S_s6_213), .c_out(C_s6_213));
FA FA_s6_214(.A(comb[15][6]), .B(comb[16][5]), .c_in(comb[17][4]), .S(S_s6_214), .c_out(C_s6_214));
FA FA_s6_215(.A(comb[18][3]), .B(comb[19][2]), .c_in(comb[20][1]), .S(S_s6_215), .c_out(C_s6_215));
FA FA_s6_220(.A(S_s7_223), .B(S_s7_222), .c_in(S_s7_221), .S(S_s6_220), .c_out(C_s6_220));
FA FA_s6_221(.A(S_s7_220), .B(C_s7_212), .c_in(C_s7_211), .S(S_s6_221), .c_out(C_s6_221));
FA FA_s6_222(.A(C_s7_210), .B(comb[11][11]), .c_in(comb[12][10]), .S(S_s6_222), .c_out(C_s6_222));
FA FA_s6_223(.A(comb[13][9]), .B(comb[14][8]), .c_in(comb[15][7]), .S(S_s6_223), .c_out(C_s6_223));
FA FA_s6_224(.A(comb[16][6]), .B(comb[17][5]), .c_in(comb[18][4]), .S(S_s6_224), .c_out(C_s6_224));
FA FA_s6_225(.A(comb[19][3]), .B(comb[20][2]), .c_in(comb[21][1]), .S(S_s6_225), .c_out(C_s6_225));
FA FA_s6_230(.A(S_s7_234), .B(S_s7_233), .c_in(S_s7_232), .S(S_s6_230), .c_out(C_s6_230));
FA FA_s6_231(.A(S_s7_231), .B(S_s7_230), .c_in(C_s7_223), .S(S_s6_231), .c_out(C_s6_231));
FA FA_s6_232(.A(C_s7_222), .B(C_s7_221), .c_in(C_s7_220), .S(S_s6_232), .c_out(C_s6_232));
FA FA_s6_233(.A(comb[14][9]), .B(comb[15][8]), .c_in(comb[16][7]), .S(S_s6_233), .c_out(C_s6_233));
FA FA_s6_234(.A(comb[17][6]), .B(comb[18][5]), .c_in(comb[19][4]), .S(S_s6_234), .c_out(C_s6_234));
FA FA_s6_235(.A(comb[20][3]), .B(comb[21][2]), .c_in(comb[22][1]), .S(S_s6_235), .c_out(C_s6_235));
FA FA_s6_240(.A(S_s7_245), .B(S_s7_244), .c_in(S_s7_243), .S(S_s6_240), .c_out(C_s6_240));
FA FA_s6_241(.A(S_s7_242), .B(S_s7_241), .c_in(S_s7_240), .S(S_s6_241), .c_out(C_s6_241));
FA FA_s6_242(.A(C_s7_234), .B(C_s7_233), .c_in(C_s7_232), .S(S_s6_242), .c_out(C_s6_242));
FA FA_s6_243(.A(C_s7_231), .B(C_s7_230), .c_in(comb[17][7]), .S(S_s6_243), .c_out(C_s6_243));
FA FA_s6_244(.A(comb[18][6]), .B(comb[19][5]), .c_in(comb[20][4]), .S(S_s6_244), .c_out(C_s6_244));
FA FA_s6_245(.A(comb[21][3]), .B(comb[22][2]), .c_in(comb[23][1]), .S(S_s6_245), .c_out(C_s6_245));
FA FA_s6_250(.A(S_s7_256), .B(S_s7_255), .c_in(S_s7_254), .S(S_s6_250), .c_out(C_s6_250));
FA FA_s6_251(.A(S_s7_253), .B(S_s7_252), .c_in(S_s7_251), .S(S_s6_251), .c_out(C_s6_251));
FA FA_s6_252(.A(S_s7_250), .B(C_s7_245), .c_in(C_s7_244), .S(S_s6_252), .c_out(C_s6_252));
FA FA_s6_253(.A(C_s7_243), .B(C_s7_242), .c_in(C_s7_241), .S(S_s6_253), .c_out(C_s6_253));
FA FA_s6_254(.A(C_s7_240), .B(comb[20][5]), .c_in(comb[21][4]), .S(S_s6_254), .c_out(C_s6_254));
FA FA_s6_255(.A(comb[22][3]), .B(comb[23][2]), .c_in(comb[24][1]), .S(S_s6_255), .c_out(C_s6_255));
FA FA_s6_260(.A(S_s7_267), .B(S_s7_266), .c_in(S_s7_265), .S(S_s6_260), .c_out(C_s6_260));
FA FA_s6_261(.A(S_s7_264), .B(S_s7_263), .c_in(S_s7_262), .S(S_s6_261), .c_out(C_s6_261));
FA FA_s6_262(.A(S_s7_261), .B(S_s7_260), .c_in(C_s7_256), .S(S_s6_262), .c_out(C_s6_262));
FA FA_s6_263(.A(C_s7_255), .B(C_s7_254), .c_in(C_s7_253), .S(S_s6_263), .c_out(C_s6_263));
FA FA_s6_264(.A(C_s7_252), .B(C_s7_251), .c_in(C_s7_250), .S(S_s6_264), .c_out(C_s6_264));
FA FA_s6_265(.A(comb[23][3]), .B(comb[24][2]), .c_in(comb[25][1]), .S(S_s6_265), .c_out(C_s6_265));
FA FA_s6_270(.A(S_s7_278), .B(S_s7_277), .c_in(S_s7_276), .S(S_s6_270), .c_out(C_s6_270));
FA FA_s6_271(.A(S_s7_275), .B(S_s7_274), .c_in(S_s7_273), .S(S_s6_271), .c_out(C_s6_271));
FA FA_s6_272(.A(S_s7_272), .B(S_s7_271), .c_in(S_s7_270), .S(S_s6_272), .c_out(C_s6_272));
FA FA_s6_273(.A(C_s7_267), .B(C_s7_266), .c_in(C_s7_265), .S(S_s6_273), .c_out(C_s6_273));
FA FA_s6_274(.A(C_s7_264), .B(C_s7_263), .c_in(C_s7_262), .S(S_s6_274), .c_out(C_s6_274));
FA FA_s6_275(.A(C_s7_261), .B(C_s7_260), .c_in(comb[26][1]), .S(S_s6_275), .c_out(C_s6_275));
FA FA_s6_280(.A(S_s7_288), .B(S_s7_287), .c_in(S_s7_286), .S(S_s6_280), .c_out(C_s6_280));
FA FA_s6_281(.A(S_s7_285), .B(S_s7_284), .c_in(S_s7_283), .S(S_s6_281), .c_out(C_s6_281));
FA FA_s6_282(.A(S_s7_282), .B(S_s7_281), .c_in(S_s7_280), .S(S_s6_282), .c_out(C_s6_282));
FA FA_s6_283(.A(C_s7_278), .B(C_s7_277), .c_in(C_s7_276), .S(S_s6_283), .c_out(C_s6_283));
FA FA_s6_284(.A(C_s7_275), .B(C_s7_274), .c_in(C_s7_273), .S(S_s6_284), .c_out(C_s6_284));
FA FA_s6_285(.A(C_s7_272), .B(C_s7_271), .c_in(C_s7_270), .S(S_s6_285), .c_out(C_s6_285));
FA FA_s6_290(.A(S_s7_298), .B(S_s7_297), .c_in(S_s7_296), .S(S_s6_290), .c_out(C_s6_290));
FA FA_s6_291(.A(S_s7_295), .B(S_s7_294), .c_in(S_s7_293), .S(S_s6_291), .c_out(C_s6_291));
FA FA_s6_292(.A(S_s7_292), .B(S_s7_291), .c_in(S_s7_290), .S(S_s6_292), .c_out(C_s6_292));
FA FA_s6_293(.A(C_s7_288), .B(C_s7_287), .c_in(C_s7_286), .S(S_s6_293), .c_out(C_s6_293));
FA FA_s6_294(.A(C_s7_285), .B(C_s7_284), .c_in(C_s7_283), .S(S_s6_294), .c_out(C_s6_294));
FA FA_s6_295(.A(C_s7_282), .B(C_s7_281), .c_in(C_s7_280), .S(S_s6_295), .c_out(C_s6_295));
FA FA_s6_300(.A(S_s7_308), .B(S_s7_307), .c_in(S_s7_306), .S(S_s6_300), .c_out(C_s6_300));
FA FA_s6_301(.A(S_s7_305), .B(S_s7_304), .c_in(S_s7_303), .S(S_s6_301), .c_out(C_s6_301));
FA FA_s6_302(.A(S_s7_302), .B(S_s7_301), .c_in(S_s7_300), .S(S_s6_302), .c_out(C_s6_302));
FA FA_s6_303(.A(C_s7_298), .B(C_s7_297), .c_in(C_s7_296), .S(S_s6_303), .c_out(C_s6_303));
FA FA_s6_304(.A(C_s7_295), .B(C_s7_294), .c_in(C_s7_293), .S(S_s6_304), .c_out(C_s6_304));
FA FA_s6_305(.A(C_s7_292), .B(C_s7_291), .c_in(C_s7_290), .S(S_s6_305), .c_out(C_s6_305));
FA FA_s6_310(.A(S_s7_318), .B(S_s7_317), .c_in(S_s7_316), .S(S_s6_310), .c_out(C_s6_310));
FA FA_s6_311(.A(S_s7_315), .B(S_s7_314), .c_in(S_s7_313), .S(S_s6_311), .c_out(C_s6_311));
FA FA_s6_312(.A(S_s7_312), .B(S_s7_311), .c_in(S_s7_310), .S(S_s6_312), .c_out(C_s6_312));
FA FA_s6_313(.A(C_s7_308), .B(C_s7_307), .c_in(C_s7_306), .S(S_s6_313), .c_out(C_s6_313));
FA FA_s6_314(.A(C_s7_305), .B(C_s7_304), .c_in(C_s7_303), .S(S_s6_314), .c_out(C_s6_314));
FA FA_s6_315(.A(C_s7_302), .B(C_s7_301), .c_in(C_s7_300), .S(S_s6_315), .c_out(C_s6_315));
FA FA_s6_320(.A(S_s7_328), .B(S_s7_327), .c_in(S_s7_326), .S(S_s6_320), .c_out(C_s6_320));
FA FA_s6_321(.A(S_s7_325), .B(S_s7_324), .c_in(S_s7_323), .S(S_s6_321), .c_out(C_s6_321));
FA FA_s6_322(.A(S_s7_322), .B(S_s7_321), .c_in(S_s7_320), .S(S_s6_322), .c_out(C_s6_322));
FA FA_s6_323(.A(C_s7_318), .B(C_s7_317), .c_in(C_s7_316), .S(S_s6_323), .c_out(C_s6_323));
FA FA_s6_324(.A(C_s7_315), .B(C_s7_314), .c_in(C_s7_313), .S(S_s6_324), .c_out(C_s6_324));
FA FA_s6_325(.A(C_s7_312), .B(C_s7_311), .c_in(C_s7_310), .S(S_s6_325), .c_out(C_s6_325));
FA FA_s6_330(.A(S_s7_338), .B(S_s7_337), .c_in(S_s7_336), .S(S_s6_330), .c_out(C_s6_330));
FA FA_s6_331(.A(S_s7_335), .B(S_s7_334), .c_in(S_s7_333), .S(S_s6_331), .c_out(C_s6_331));
FA FA_s6_332(.A(S_s7_332), .B(S_s7_331), .c_in(S_s7_330), .S(S_s6_332), .c_out(C_s6_332));
FA FA_s6_333(.A(C_s7_328), .B(C_s7_327), .c_in(C_s7_326), .S(S_s6_333), .c_out(C_s6_333));
FA FA_s6_334(.A(C_s7_325), .B(C_s7_324), .c_in(C_s7_323), .S(S_s6_334), .c_out(C_s6_334));
FA FA_s6_335(.A(C_s7_322), .B(C_s7_321), .c_in(C_s7_320), .S(S_s6_335), .c_out(C_s6_335));
FA FA_s6_340(.A(S_s7_348), .B(S_s7_347), .c_in(S_s7_346), .S(S_s6_340), .c_out(C_s6_340));
FA FA_s6_341(.A(S_s7_345), .B(S_s7_344), .c_in(S_s7_343), .S(S_s6_341), .c_out(C_s6_341));
FA FA_s6_342(.A(S_s7_342), .B(S_s7_341), .c_in(S_s7_340), .S(S_s6_342), .c_out(C_s6_342));
FA FA_s6_343(.A(C_s7_338), .B(C_s7_337), .c_in(C_s7_336), .S(S_s6_343), .c_out(C_s6_343));
FA FA_s6_344(.A(C_s7_335), .B(C_s7_334), .c_in(C_s7_333), .S(S_s6_344), .c_out(C_s6_344));
FA FA_s6_345(.A(C_s7_332), .B(C_s7_331), .c_in(C_s7_330), .S(S_s6_345), .c_out(C_s6_345));
FA FA_s6_350(.A(S_s7_358), .B(S_s7_357), .c_in(S_s7_356), .S(S_s6_350), .c_out(C_s6_350));
FA FA_s6_351(.A(S_s7_355), .B(S_s7_354), .c_in(S_s7_353), .S(S_s6_351), .c_out(C_s6_351));
FA FA_s6_352(.A(S_s7_352), .B(S_s7_351), .c_in(S_s7_350), .S(S_s6_352), .c_out(C_s6_352));
FA FA_s6_353(.A(C_s7_348), .B(C_s7_347), .c_in(C_s7_346), .S(S_s6_353), .c_out(C_s6_353));
FA FA_s6_354(.A(C_s7_345), .B(C_s7_344), .c_in(C_s7_343), .S(S_s6_354), .c_out(C_s6_354));
FA FA_s6_355(.A(C_s7_342), .B(C_s7_341), .c_in(C_s7_340), .S(S_s6_355), .c_out(C_s6_355));
FA FA_s6_360(.A(S_s7_368), .B(S_s7_367), .c_in(S_s7_366), .S(S_s6_360), .c_out(C_s6_360));
FA FA_s6_361(.A(S_s7_365), .B(S_s7_364), .c_in(S_s7_363), .S(S_s6_361), .c_out(C_s6_361));
FA FA_s6_362(.A(S_s7_362), .B(S_s7_361), .c_in(S_s7_360), .S(S_s6_362), .c_out(C_s6_362));
FA FA_s6_363(.A(C_s7_358), .B(C_s7_357), .c_in(C_s7_356), .S(S_s6_363), .c_out(C_s6_363));
FA FA_s6_364(.A(C_s7_355), .B(C_s7_354), .c_in(C_s7_353), .S(S_s6_364), .c_out(C_s6_364));
FA FA_s6_365(.A(C_s7_352), .B(C_s7_351), .c_in(C_s7_350), .S(S_s6_365), .c_out(C_s6_365));
FA FA_s6_370(.A(S_s7_377), .B(S_s7_376), .c_in(S_s7_375), .S(S_s6_370), .c_out(C_s6_370));
FA FA_s6_371(.A(S_s7_374), .B(S_s7_373), .c_in(S_s7_372), .S(S_s6_371), .c_out(C_s6_371));
FA FA_s6_372(.A(S_s7_371), .B(S_s7_370), .c_in(C_s7_368), .S(S_s6_372), .c_out(C_s6_372));
FA FA_s6_373(.A(C_s7_367), .B(C_s7_366), .c_in(C_s7_365), .S(S_s6_373), .c_out(C_s6_373));
FA FA_s6_374(.A(C_s7_364), .B(C_s7_363), .c_in(C_s7_362), .S(S_s6_374), .c_out(C_s6_374));
FA FA_s6_375(.A(C_s7_361), .B(C_s7_360), .c_in(comb[30][7]), .S(S_s6_375), .c_out(C_s6_375));
FA FA_s6_380(.A(S_s7_386), .B(S_s7_385), .c_in(S_s7_384), .S(S_s6_380), .c_out(C_s6_380));
FA FA_s6_381(.A(S_s7_383), .B(S_s7_382), .c_in(S_s7_381), .S(S_s6_381), .c_out(C_s6_381));
FA FA_s6_382(.A(S_s7_380), .B(C_s7_377), .c_in(C_s7_376), .S(S_s6_382), .c_out(C_s6_382));
FA FA_s6_383(.A(C_s7_375), .B(C_s7_374), .c_in(C_s7_373), .S(S_s6_383), .c_out(C_s6_383));
FA FA_s6_384(.A(C_s7_372), .B(C_s7_371), .c_in(C_s7_370), .S(S_s6_384), .c_out(C_s6_384));
FA FA_s6_385(.A(comb[28][10]), .B(comb[29][9]), .c_in(comb[30][8]), .S(S_s6_385), .c_out(C_s6_385));
FA FA_s6_390(.A(S_s7_395), .B(S_s7_394), .c_in(S_s7_393), .S(S_s6_390), .c_out(C_s6_390));
FA FA_s6_391(.A(S_s7_392), .B(S_s7_391), .c_in(S_s7_390), .S(S_s6_391), .c_out(C_s6_391));
FA FA_s6_392(.A(C_s7_386), .B(C_s7_385), .c_in(C_s7_384), .S(S_s6_392), .c_out(C_s6_392));
FA FA_s6_393(.A(C_s7_383), .B(C_s7_382), .c_in(C_s7_381), .S(S_s6_393), .c_out(C_s6_393));
FA FA_s6_394(.A(C_s7_380), .B(comb[26][13]), .c_in(comb[27][12]), .S(S_s6_394), .c_out(C_s6_394));
FA FA_s6_395(.A(comb[28][11]), .B(comb[29][10]), .c_in(comb[30][9]), .S(S_s6_395), .c_out(C_s6_395));
FA FA_s6_400(.A(S_s7_404), .B(S_s7_403), .c_in(S_s7_402), .S(S_s6_400), .c_out(C_s6_400));
FA FA_s6_401(.A(S_s7_401), .B(S_s7_400), .c_in(C_s7_395), .S(S_s6_401), .c_out(C_s6_401));
FA FA_s6_402(.A(C_s7_394), .B(C_s7_393), .c_in(C_s7_392), .S(S_s6_402), .c_out(C_s6_402));
FA FA_s6_403(.A(C_s7_391), .B(C_s7_390), .c_in(comb[24][16]), .S(S_s6_403), .c_out(C_s6_403));
FA FA_s6_404(.A(comb[25][15]), .B(comb[26][14]), .c_in(comb[27][13]), .S(S_s6_404), .c_out(C_s6_404));
FA FA_s6_405(.A(comb[28][12]), .B(comb[29][11]), .c_in(comb[30][10]), .S(S_s6_405), .c_out(C_s6_405));
FA FA_s6_410(.A(S_s7_413), .B(S_s7_412), .c_in(S_s7_411), .S(S_s6_410), .c_out(C_s6_410));
FA FA_s6_411(.A(S_s7_410), .B(C_s7_404), .c_in(C_s7_403), .S(S_s6_411), .c_out(C_s6_411));
FA FA_s6_412(.A(C_s7_402), .B(C_s7_401), .c_in(C_s7_400), .S(S_s6_412), .c_out(C_s6_412));
FA FA_s6_413(.A(comb[22][19]), .B(comb[23][18]), .c_in(comb[24][17]), .S(S_s6_413), .c_out(C_s6_413));
FA FA_s6_414(.A(comb[25][16]), .B(comb[26][15]), .c_in(comb[27][14]), .S(S_s6_414), .c_out(C_s6_414));
FA FA_s6_415(.A(comb[28][13]), .B(comb[29][12]), .c_in(comb[30][11]), .S(S_s6_415), .c_out(C_s6_415));
FA FA_s6_420(.A(S_s7_422), .B(S_s7_421), .c_in(S_s7_420), .S(S_s6_420), .c_out(C_s6_420));
FA FA_s6_421(.A(C_s7_413), .B(C_s7_412), .c_in(C_s7_411), .S(S_s6_421), .c_out(C_s6_421));
FA FA_s6_422(.A(C_s7_410), .B(comb[20][22]), .c_in(comb[21][21]), .S(S_s6_422), .c_out(C_s6_422));
FA FA_s6_423(.A(comb[22][20]), .B(comb[23][19]), .c_in(comb[24][18]), .S(S_s6_423), .c_out(C_s6_423));
FA FA_s6_424(.A(comb[25][17]), .B(comb[26][16]), .c_in(comb[27][15]), .S(S_s6_424), .c_out(C_s6_424));
FA FA_s6_425(.A(comb[28][14]), .B(comb[29][13]), .c_in(comb[30][12]), .S(S_s6_425), .c_out(C_s6_425));
FA FA_s6_430(.A(S_s7_431), .B(S_s7_430), .c_in(C_s7_422), .S(S_s6_430), .c_out(C_s6_430));
FA FA_s6_431(.A(C_s7_421), .B(C_s7_420), .c_in(comb[18][25]), .S(S_s6_431), .c_out(C_s6_431));
FA FA_s6_432(.A(comb[19][24]), .B(comb[20][23]), .c_in(comb[21][22]), .S(S_s6_432), .c_out(C_s6_432));
FA FA_s6_433(.A(comb[22][21]), .B(comb[23][20]), .c_in(comb[24][19]), .S(S_s6_433), .c_out(C_s6_433));
FA FA_s6_434(.A(comb[25][18]), .B(comb[26][17]), .c_in(comb[27][16]), .S(S_s6_434), .c_out(C_s6_434));
FA FA_s6_435(.A(comb[28][15]), .B(comb[29][14]), .c_in(comb[30][13]), .S(S_s6_435), .c_out(C_s6_435));
FA FA_s6_440(.A(S_s7_440), .B(C_s7_431), .c_in(C_s7_430), .S(S_s6_440), .c_out(C_s6_440));
FA FA_s6_441(.A(comb[16][28]), .B(comb[17][27]), .c_in(comb[18][26]), .S(S_s6_441), .c_out(C_s6_441));
FA FA_s6_442(.A(comb[19][25]), .B(comb[20][24]), .c_in(comb[21][23]), .S(S_s6_442), .c_out(C_s6_442));
FA FA_s6_443(.A(comb[22][22]), .B(comb[23][21]), .c_in(comb[24][20]), .S(S_s6_443), .c_out(C_s6_443));
FA FA_s6_444(.A(comb[25][19]), .B(comb[26][18]), .c_in(comb[27][17]), .S(S_s6_444), .c_out(C_s6_444));
FA FA_s6_445(.A(comb[28][16]), .B(comb[29][15]), .c_in(comb[30][14]), .S(S_s6_445), .c_out(C_s6_445));
FA FA_s6_450(.A(C_s7_440), .B(comb[14][31]), .c_in(comb[15][30]), .S(S_s6_450), .c_out(C_s6_450));
FA FA_s6_451(.A(comb[16][29]), .B(comb[17][28]), .c_in(comb[18][27]), .S(S_s6_451), .c_out(C_s6_451));
FA FA_s6_452(.A(comb[19][26]), .B(comb[20][25]), .c_in(comb[21][24]), .S(S_s6_452), .c_out(C_s6_452));
FA FA_s6_453(.A(comb[22][23]), .B(comb[23][22]), .c_in(comb[24][21]), .S(S_s6_453), .c_out(C_s6_453));
FA FA_s6_454(.A(comb[25][20]), .B(comb[26][19]), .c_in(comb[27][18]), .S(S_s6_454), .c_out(C_s6_454));
FA FA_s6_455(.A(comb[28][17]), .B(comb[29][16]), .c_in(comb[30][15]), .S(S_s6_455), .c_out(C_s6_455));
FA FA_s6_460(.A(comb[15][31]), .B(comb[16][30]), .c_in(comb[17][29]), .S(S_s6_460), .c_out(C_s6_460));
FA FA_s6_461(.A(comb[18][28]), .B(comb[19][27]), .c_in(comb[20][26]), .S(S_s6_461), .c_out(C_s6_461));
FA FA_s6_462(.A(comb[21][25]), .B(comb[22][24]), .c_in(comb[23][23]), .S(S_s6_462), .c_out(C_s6_462));
FA FA_s6_463(.A(comb[24][22]), .B(comb[25][21]), .c_in(comb[26][20]), .S(S_s6_463), .c_out(C_s6_463));
FA FA_s6_464(.A(comb[27][19]), .B(comb[28][18]), .c_in(comb[29][17]), .S(S_s6_464), .c_out(C_s6_464));
FA FA_s6_470(.A(comb[16][31]), .B(comb[17][30]), .c_in(comb[18][29]), .S(S_s6_470), .c_out(C_s6_470));
FA FA_s6_471(.A(comb[19][28]), .B(comb[20][27]), .c_in(comb[21][26]), .S(S_s6_471), .c_out(C_s6_471));
FA FA_s6_472(.A(comb[22][25]), .B(comb[23][24]), .c_in(comb[24][23]), .S(S_s6_472), .c_out(C_s6_472));
FA FA_s6_473(.A(comb[25][22]), .B(comb[26][21]), .c_in(comb[27][20]), .S(S_s6_473), .c_out(C_s6_473));
FA FA_s6_480(.A(comb[17][31]), .B(comb[18][30]), .c_in(comb[19][29]), .S(S_s6_480), .c_out(C_s6_480));
FA FA_s6_481(.A(comb[20][28]), .B(comb[21][27]), .c_in(comb[22][26]), .S(S_s6_481), .c_out(C_s6_481));
FA FA_s6_482(.A(comb[23][25]), .B(comb[24][24]), .c_in(comb[25][23]), .S(S_s6_482), .c_out(C_s6_482));
FA FA_s6_490(.A(comb[18][31]), .B(comb[19][30]), .c_in(comb[20][29]), .S(S_s6_490), .c_out(C_s6_490));
FA FA_s6_491(.A(comb[21][28]), .B(comb[22][27]), .c_in(comb[23][26]), .S(S_s6_491), .c_out(C_s6_491));
FA FA_s6_500(.A(comb[19][31]), .B(comb[20][30]), .c_in(comb[21][29]), .S(S_s6_500), .c_out(C_s6_500));
// stage 6 end ======================================================================= 

// stage 5 begin ======================================================================= 
HA HA_s5_90(.A(comb[0][9]), .B(comb[1][8]), .S(S_s5_90), .c_out(C_s5_90));
FA FA_s5_100(.A(comb[0][10]), .B(comb[1][9]), .c_in(comb[2][8]), .S(S_s5_100), .c_out(C_s5_100));
HA HA_s5_101(.A(comb[3][7]), .B(comb[4][6]), .S(S_s5_101), .c_out(C_s5_101));
FA FA_s5_110(.A(comb[0][11]), .B(comb[1][10]), .c_in(comb[2][9]), .S(S_s5_110), .c_out(C_s5_110));
FA FA_s5_111(.A(comb[3][8]), .B(comb[4][7]), .c_in(comb[5][6]), .S(S_s5_111), .c_out(C_s5_111));
HA HA_s5_112(.A(comb[6][5]), .B(comb[7][4]), .S(S_s5_112), .c_out(C_s5_112));
FA FA_s5_120(.A(comb[0][12]), .B(comb[1][11]), .c_in(comb[2][10]), .S(S_s5_120), .c_out(C_s5_120));
FA FA_s5_121(.A(comb[3][9]), .B(comb[4][8]), .c_in(comb[5][7]), .S(S_s5_121), .c_out(C_s5_121));
FA FA_s5_122(.A(comb[6][6]), .B(comb[7][5]), .c_in(comb[8][4]), .S(S_s5_122), .c_out(C_s5_122));
HA HA_s5_123(.A(comb[9][3]), .B(comb[10][2]), .S(S_s5_123), .c_out(C_s5_123));
FA FA_s5_130(.A(S_s6_130), .B(comb[2][11]), .c_in(comb[3][10]), .S(S_s5_130), .c_out(C_s5_130));
FA FA_s5_131(.A(comb[4][9]), .B(comb[5][8]), .c_in(comb[6][7]), .S(S_s5_131), .c_out(C_s5_131));
FA FA_s5_132(.A(comb[7][6]), .B(comb[8][5]), .c_in(comb[9][4]), .S(S_s5_132), .c_out(C_s5_132));
FA FA_s5_133(.A(comb[10][3]), .B(comb[11][2]), .c_in(comb[12][1]), .S(S_s5_133), .c_out(C_s5_133));
FA FA_s5_140(.A(S_s6_141), .B(S_s6_140), .c_in(C_s6_130), .S(S_s5_140), .c_out(C_s5_140));
FA FA_s5_141(.A(comb[5][9]), .B(comb[6][8]), .c_in(comb[7][7]), .S(S_s5_141), .c_out(C_s5_141));
FA FA_s5_142(.A(comb[8][6]), .B(comb[9][5]), .c_in(comb[10][4]), .S(S_s5_142), .c_out(C_s5_142));
FA FA_s5_143(.A(comb[11][3]), .B(comb[12][2]), .c_in(comb[13][1]), .S(S_s5_143), .c_out(C_s5_143));
FA FA_s5_150(.A(S_s6_152), .B(S_s6_151), .c_in(S_s6_150), .S(S_s5_150), .c_out(C_s5_150));
FA FA_s5_151(.A(C_s6_141), .B(C_s6_140), .c_in(comb[8][7]), .S(S_s5_151), .c_out(C_s5_151));
FA FA_s5_152(.A(comb[9][6]), .B(comb[10][5]), .c_in(comb[11][4]), .S(S_s5_152), .c_out(C_s5_152));
FA FA_s5_153(.A(comb[12][3]), .B(comb[13][2]), .c_in(comb[14][1]), .S(S_s5_153), .c_out(C_s5_153));
FA FA_s5_160(.A(S_s6_163), .B(S_s6_162), .c_in(S_s6_161), .S(S_s5_160), .c_out(C_s5_160));
FA FA_s5_161(.A(S_s6_160), .B(C_s6_152), .c_in(C_s6_151), .S(S_s5_161), .c_out(C_s5_161));
FA FA_s5_162(.A(C_s6_150), .B(comb[11][5]), .c_in(comb[12][4]), .S(S_s5_162), .c_out(C_s5_162));
FA FA_s5_163(.A(comb[13][3]), .B(comb[14][2]), .c_in(comb[15][1]), .S(S_s5_163), .c_out(C_s5_163));
FA FA_s5_170(.A(S_s6_174), .B(S_s6_173), .c_in(S_s6_172), .S(S_s5_170), .c_out(C_s5_170));
FA FA_s5_171(.A(S_s6_171), .B(S_s6_170), .c_in(C_s6_163), .S(S_s5_171), .c_out(C_s5_171));
FA FA_s5_172(.A(C_s6_162), .B(C_s6_161), .c_in(C_s6_160), .S(S_s5_172), .c_out(C_s5_172));
FA FA_s5_173(.A(comb[14][3]), .B(comb[15][2]), .c_in(comb[16][1]), .S(S_s5_173), .c_out(C_s5_173));
FA FA_s5_180(.A(S_s6_185), .B(S_s6_184), .c_in(S_s6_183), .S(S_s5_180), .c_out(C_s5_180));
FA FA_s5_181(.A(S_s6_182), .B(S_s6_181), .c_in(S_s6_180), .S(S_s5_181), .c_out(C_s5_181));
FA FA_s5_182(.A(C_s6_174), .B(C_s6_173), .c_in(C_s6_172), .S(S_s5_182), .c_out(C_s5_182));
FA FA_s5_183(.A(C_s6_171), .B(C_s6_170), .c_in(comb[17][1]), .S(S_s5_183), .c_out(C_s5_183));
FA FA_s5_190(.A(S_s6_195), .B(S_s6_194), .c_in(S_s6_193), .S(S_s5_190), .c_out(C_s5_190));
FA FA_s5_191(.A(S_s6_192), .B(S_s6_191), .c_in(S_s6_190), .S(S_s5_191), .c_out(C_s5_191));
FA FA_s5_192(.A(C_s6_185), .B(C_s6_184), .c_in(C_s6_183), .S(S_s5_192), .c_out(C_s5_192));
FA FA_s5_193(.A(C_s6_182), .B(C_s6_181), .c_in(C_s6_180), .S(S_s5_193), .c_out(C_s5_193));
FA FA_s5_200(.A(S_s6_205), .B(S_s6_204), .c_in(S_s6_203), .S(S_s5_200), .c_out(C_s5_200));
FA FA_s5_201(.A(S_s6_202), .B(S_s6_201), .c_in(S_s6_200), .S(S_s5_201), .c_out(C_s5_201));
FA FA_s5_202(.A(C_s6_195), .B(C_s6_194), .c_in(C_s6_193), .S(S_s5_202), .c_out(C_s5_202));
FA FA_s5_203(.A(C_s6_192), .B(C_s6_191), .c_in(C_s6_190), .S(S_s5_203), .c_out(C_s5_203));
FA FA_s5_210(.A(S_s6_215), .B(S_s6_214), .c_in(S_s6_213), .S(S_s5_210), .c_out(C_s5_210));
FA FA_s5_211(.A(S_s6_212), .B(S_s6_211), .c_in(S_s6_210), .S(S_s5_211), .c_out(C_s5_211));
FA FA_s5_212(.A(C_s6_205), .B(C_s6_204), .c_in(C_s6_203), .S(S_s5_212), .c_out(C_s5_212));
FA FA_s5_213(.A(C_s6_202), .B(C_s6_201), .c_in(C_s6_200), .S(S_s5_213), .c_out(C_s5_213));
FA FA_s5_220(.A(S_s6_225), .B(S_s6_224), .c_in(S_s6_223), .S(S_s5_220), .c_out(C_s5_220));
FA FA_s5_221(.A(S_s6_222), .B(S_s6_221), .c_in(S_s6_220), .S(S_s5_221), .c_out(C_s5_221));
FA FA_s5_222(.A(C_s6_215), .B(C_s6_214), .c_in(C_s6_213), .S(S_s5_222), .c_out(C_s5_222));
FA FA_s5_223(.A(C_s6_212), .B(C_s6_211), .c_in(C_s6_210), .S(S_s5_223), .c_out(C_s5_223));
FA FA_s5_230(.A(S_s6_235), .B(S_s6_234), .c_in(S_s6_233), .S(S_s5_230), .c_out(C_s5_230));
FA FA_s5_231(.A(S_s6_232), .B(S_s6_231), .c_in(S_s6_230), .S(S_s5_231), .c_out(C_s5_231));
FA FA_s5_232(.A(C_s6_225), .B(C_s6_224), .c_in(C_s6_223), .S(S_s5_232), .c_out(C_s5_232));
FA FA_s5_233(.A(C_s6_222), .B(C_s6_221), .c_in(C_s6_220), .S(S_s5_233), .c_out(C_s5_233));
FA FA_s5_240(.A(S_s6_245), .B(S_s6_244), .c_in(S_s6_243), .S(S_s5_240), .c_out(C_s5_240));
FA FA_s5_241(.A(S_s6_242), .B(S_s6_241), .c_in(S_s6_240), .S(S_s5_241), .c_out(C_s5_241));
FA FA_s5_242(.A(C_s6_235), .B(C_s6_234), .c_in(C_s6_233), .S(S_s5_242), .c_out(C_s5_242));
FA FA_s5_243(.A(C_s6_232), .B(C_s6_231), .c_in(C_s6_230), .S(S_s5_243), .c_out(C_s5_243));
FA FA_s5_250(.A(S_s6_255), .B(S_s6_254), .c_in(S_s6_253), .S(S_s5_250), .c_out(C_s5_250));
FA FA_s5_251(.A(S_s6_252), .B(S_s6_251), .c_in(S_s6_250), .S(S_s5_251), .c_out(C_s5_251));
FA FA_s5_252(.A(C_s6_245), .B(C_s6_244), .c_in(C_s6_243), .S(S_s5_252), .c_out(C_s5_252));
FA FA_s5_253(.A(C_s6_242), .B(C_s6_241), .c_in(C_s6_240), .S(S_s5_253), .c_out(C_s5_253));
FA FA_s5_260(.A(S_s6_265), .B(S_s6_264), .c_in(S_s6_263), .S(S_s5_260), .c_out(C_s5_260));
FA FA_s5_261(.A(S_s6_262), .B(S_s6_261), .c_in(S_s6_260), .S(S_s5_261), .c_out(C_s5_261));
FA FA_s5_262(.A(C_s6_255), .B(C_s6_254), .c_in(C_s6_253), .S(S_s5_262), .c_out(C_s5_262));
FA FA_s5_263(.A(C_s6_252), .B(C_s6_251), .c_in(C_s6_250), .S(S_s5_263), .c_out(C_s5_263));
FA FA_s5_270(.A(S_s6_275), .B(S_s6_274), .c_in(S_s6_273), .S(S_s5_270), .c_out(C_s5_270));
FA FA_s5_271(.A(S_s6_272), .B(S_s6_271), .c_in(S_s6_270), .S(S_s5_271), .c_out(C_s5_271));
FA FA_s5_272(.A(C_s6_265), .B(C_s6_264), .c_in(C_s6_263), .S(S_s5_272), .c_out(C_s5_272));
FA FA_s5_273(.A(C_s6_262), .B(C_s6_261), .c_in(C_s6_260), .S(S_s5_273), .c_out(C_s5_273));
FA FA_s5_280(.A(S_s6_285), .B(S_s6_284), .c_in(S_s6_283), .S(S_s5_280), .c_out(C_s5_280));
FA FA_s5_281(.A(S_s6_282), .B(S_s6_281), .c_in(S_s6_280), .S(S_s5_281), .c_out(C_s5_281));
FA FA_s5_282(.A(C_s6_275), .B(C_s6_274), .c_in(C_s6_273), .S(S_s5_282), .c_out(C_s5_282));
FA FA_s5_283(.A(C_s6_272), .B(C_s6_271), .c_in(C_s6_270), .S(S_s5_283), .c_out(C_s5_283));
FA FA_s5_290(.A(S_s6_295), .B(S_s6_294), .c_in(S_s6_293), .S(S_s5_290), .c_out(C_s5_290));
FA FA_s5_291(.A(S_s6_292), .B(S_s6_291), .c_in(S_s6_290), .S(S_s5_291), .c_out(C_s5_291));
FA FA_s5_292(.A(C_s6_285), .B(C_s6_284), .c_in(C_s6_283), .S(S_s5_292), .c_out(C_s5_292));
FA FA_s5_293(.A(C_s6_282), .B(C_s6_281), .c_in(C_s6_280), .S(S_s5_293), .c_out(C_s5_293));
FA FA_s5_300(.A(S_s6_305), .B(S_s6_304), .c_in(S_s6_303), .S(S_s5_300), .c_out(C_s5_300));
FA FA_s5_301(.A(S_s6_302), .B(S_s6_301), .c_in(S_s6_300), .S(S_s5_301), .c_out(C_s5_301));
FA FA_s5_302(.A(C_s6_295), .B(C_s6_294), .c_in(C_s6_293), .S(S_s5_302), .c_out(C_s5_302));
FA FA_s5_303(.A(C_s6_292), .B(C_s6_291), .c_in(C_s6_290), .S(S_s5_303), .c_out(C_s5_303));
FA FA_s5_310(.A(S_s6_315), .B(S_s6_314), .c_in(S_s6_313), .S(S_s5_310), .c_out(C_s5_310));
FA FA_s5_311(.A(S_s6_312), .B(S_s6_311), .c_in(S_s6_310), .S(S_s5_311), .c_out(C_s5_311));
FA FA_s5_312(.A(C_s6_305), .B(C_s6_304), .c_in(C_s6_303), .S(S_s5_312), .c_out(C_s5_312));
FA FA_s5_313(.A(C_s6_302), .B(C_s6_301), .c_in(C_s6_300), .S(S_s5_313), .c_out(C_s5_313));
FA FA_s5_320(.A(S_s6_325), .B(S_s6_324), .c_in(S_s6_323), .S(S_s5_320), .c_out(C_s5_320));
FA FA_s5_321(.A(S_s6_322), .B(S_s6_321), .c_in(S_s6_320), .S(S_s5_321), .c_out(C_s5_321));
FA FA_s5_322(.A(C_s6_315), .B(C_s6_314), .c_in(C_s6_313), .S(S_s5_322), .c_out(C_s5_322));
FA FA_s5_323(.A(C_s6_312), .B(C_s6_311), .c_in(C_s6_310), .S(S_s5_323), .c_out(C_s5_323));
FA FA_s5_330(.A(S_s6_335), .B(S_s6_334), .c_in(S_s6_333), .S(S_s5_330), .c_out(C_s5_330));
FA FA_s5_331(.A(S_s6_332), .B(S_s6_331), .c_in(S_s6_330), .S(S_s5_331), .c_out(C_s5_331));
FA FA_s5_332(.A(C_s6_325), .B(C_s6_324), .c_in(C_s6_323), .S(S_s5_332), .c_out(C_s5_332));
FA FA_s5_333(.A(C_s6_322), .B(C_s6_321), .c_in(C_s6_320), .S(S_s5_333), .c_out(C_s5_333));
FA FA_s5_340(.A(S_s6_345), .B(S_s6_344), .c_in(S_s6_343), .S(S_s5_340), .c_out(C_s5_340));
FA FA_s5_341(.A(S_s6_342), .B(S_s6_341), .c_in(S_s6_340), .S(S_s5_341), .c_out(C_s5_341));
FA FA_s5_342(.A(C_s6_335), .B(C_s6_334), .c_in(C_s6_333), .S(S_s5_342), .c_out(C_s5_342));
FA FA_s5_343(.A(C_s6_332), .B(C_s6_331), .c_in(C_s6_330), .S(S_s5_343), .c_out(C_s5_343));
FA FA_s5_350(.A(S_s6_355), .B(S_s6_354), .c_in(S_s6_353), .S(S_s5_350), .c_out(C_s5_350));
FA FA_s5_351(.A(S_s6_352), .B(S_s6_351), .c_in(S_s6_350), .S(S_s5_351), .c_out(C_s5_351));
FA FA_s5_352(.A(C_s6_345), .B(C_s6_344), .c_in(C_s6_343), .S(S_s5_352), .c_out(C_s5_352));
FA FA_s5_353(.A(C_s6_342), .B(C_s6_341), .c_in(C_s6_340), .S(S_s5_353), .c_out(C_s5_353));
FA FA_s5_360(.A(S_s6_365), .B(S_s6_364), .c_in(S_s6_363), .S(S_s5_360), .c_out(C_s5_360));
FA FA_s5_361(.A(S_s6_362), .B(S_s6_361), .c_in(S_s6_360), .S(S_s5_361), .c_out(C_s5_361));
FA FA_s5_362(.A(C_s6_355), .B(C_s6_354), .c_in(C_s6_353), .S(S_s5_362), .c_out(C_s5_362));
FA FA_s5_363(.A(C_s6_352), .B(C_s6_351), .c_in(C_s6_350), .S(S_s5_363), .c_out(C_s5_363));
FA FA_s5_370(.A(S_s6_375), .B(S_s6_374), .c_in(S_s6_373), .S(S_s5_370), .c_out(C_s5_370));
FA FA_s5_371(.A(S_s6_372), .B(S_s6_371), .c_in(S_s6_370), .S(S_s5_371), .c_out(C_s5_371));
FA FA_s5_372(.A(C_s6_365), .B(C_s6_364), .c_in(C_s6_363), .S(S_s5_372), .c_out(C_s5_372));
FA FA_s5_373(.A(C_s6_362), .B(C_s6_361), .c_in(C_s6_360), .S(S_s5_373), .c_out(C_s5_373));
FA FA_s5_380(.A(S_s6_385), .B(S_s6_384), .c_in(S_s6_383), .S(S_s5_380), .c_out(C_s5_380));
FA FA_s5_381(.A(S_s6_382), .B(S_s6_381), .c_in(S_s6_380), .S(S_s5_381), .c_out(C_s5_381));
FA FA_s5_382(.A(C_s6_375), .B(C_s6_374), .c_in(C_s6_373), .S(S_s5_382), .c_out(C_s5_382));
FA FA_s5_383(.A(C_s6_372), .B(C_s6_371), .c_in(C_s6_370), .S(S_s5_383), .c_out(C_s5_383));
FA FA_s5_390(.A(S_s6_395), .B(S_s6_394), .c_in(S_s6_393), .S(S_s5_390), .c_out(C_s5_390));
FA FA_s5_391(.A(S_s6_392), .B(S_s6_391), .c_in(S_s6_390), .S(S_s5_391), .c_out(C_s5_391));
FA FA_s5_392(.A(C_s6_385), .B(C_s6_384), .c_in(C_s6_383), .S(S_s5_392), .c_out(C_s5_392));
FA FA_s5_393(.A(C_s6_382), .B(C_s6_381), .c_in(C_s6_380), .S(S_s5_393), .c_out(C_s5_393));
FA FA_s5_400(.A(S_s6_405), .B(S_s6_404), .c_in(S_s6_403), .S(S_s5_400), .c_out(C_s5_400));
FA FA_s5_401(.A(S_s6_402), .B(S_s6_401), .c_in(S_s6_400), .S(S_s5_401), .c_out(C_s5_401));
FA FA_s5_402(.A(C_s6_395), .B(C_s6_394), .c_in(C_s6_393), .S(S_s5_402), .c_out(C_s5_402));
FA FA_s5_403(.A(C_s6_392), .B(C_s6_391), .c_in(C_s6_390), .S(S_s5_403), .c_out(C_s5_403));
FA FA_s5_410(.A(S_s6_415), .B(S_s6_414), .c_in(S_s6_413), .S(S_s5_410), .c_out(C_s5_410));
FA FA_s5_411(.A(S_s6_412), .B(S_s6_411), .c_in(S_s6_410), .S(S_s5_411), .c_out(C_s5_411));
FA FA_s5_412(.A(C_s6_405), .B(C_s6_404), .c_in(C_s6_403), .S(S_s5_412), .c_out(C_s5_412));
FA FA_s5_413(.A(C_s6_402), .B(C_s6_401), .c_in(C_s6_400), .S(S_s5_413), .c_out(C_s5_413));
FA FA_s5_420(.A(S_s6_425), .B(S_s6_424), .c_in(S_s6_423), .S(S_s5_420), .c_out(C_s5_420));
FA FA_s5_421(.A(S_s6_422), .B(S_s6_421), .c_in(S_s6_420), .S(S_s5_421), .c_out(C_s5_421));
FA FA_s5_422(.A(C_s6_415), .B(C_s6_414), .c_in(C_s6_413), .S(S_s5_422), .c_out(C_s5_422));
FA FA_s5_423(.A(C_s6_412), .B(C_s6_411), .c_in(C_s6_410), .S(S_s5_423), .c_out(C_s5_423));
FA FA_s5_430(.A(S_s6_435), .B(S_s6_434), .c_in(S_s6_433), .S(S_s5_430), .c_out(C_s5_430));
FA FA_s5_431(.A(S_s6_432), .B(S_s6_431), .c_in(S_s6_430), .S(S_s5_431), .c_out(C_s5_431));
FA FA_s5_432(.A(C_s6_425), .B(C_s6_424), .c_in(C_s6_423), .S(S_s5_432), .c_out(C_s5_432));
FA FA_s5_433(.A(C_s6_422), .B(C_s6_421), .c_in(C_s6_420), .S(S_s5_433), .c_out(C_s5_433));
FA FA_s5_440(.A(S_s6_445), .B(S_s6_444), .c_in(S_s6_443), .S(S_s5_440), .c_out(C_s5_440));
FA FA_s5_441(.A(S_s6_442), .B(S_s6_441), .c_in(S_s6_440), .S(S_s5_441), .c_out(C_s5_441));
FA FA_s5_442(.A(C_s6_435), .B(C_s6_434), .c_in(C_s6_433), .S(S_s5_442), .c_out(C_s5_442));
FA FA_s5_443(.A(C_s6_432), .B(C_s6_431), .c_in(C_s6_430), .S(S_s5_443), .c_out(C_s5_443));
FA FA_s5_450(.A(S_s6_455), .B(S_s6_454), .c_in(S_s6_453), .S(S_s5_450), .c_out(C_s5_450));
FA FA_s5_451(.A(S_s6_452), .B(S_s6_451), .c_in(S_s6_450), .S(S_s5_451), .c_out(C_s5_451));
FA FA_s5_452(.A(C_s6_445), .B(C_s6_444), .c_in(C_s6_443), .S(S_s5_452), .c_out(C_s5_452));
FA FA_s5_453(.A(C_s6_442), .B(C_s6_441), .c_in(C_s6_440), .S(S_s5_453), .c_out(C_s5_453));
FA FA_s5_460(.A(S_s6_464), .B(S_s6_463), .c_in(S_s6_462), .S(S_s5_460), .c_out(C_s5_460));
FA FA_s5_461(.A(S_s6_461), .B(S_s6_460), .c_in(C_s6_455), .S(S_s5_461), .c_out(C_s5_461));
FA FA_s5_462(.A(C_s6_454), .B(C_s6_453), .c_in(C_s6_452), .S(S_s5_462), .c_out(C_s5_462));
FA FA_s5_463(.A(C_s6_451), .B(C_s6_450), .c_in(comb[30][16]), .S(S_s5_463), .c_out(C_s5_463));
FA FA_s5_470(.A(S_s6_473), .B(S_s6_472), .c_in(S_s6_471), .S(S_s5_470), .c_out(C_s5_470));
FA FA_s5_471(.A(S_s6_470), .B(C_s6_464), .c_in(C_s6_463), .S(S_s5_471), .c_out(C_s5_471));
FA FA_s5_472(.A(C_s6_462), .B(C_s6_461), .c_in(C_s6_460), .S(S_s5_472), .c_out(C_s5_472));
FA FA_s5_473(.A(comb[28][19]), .B(comb[29][18]), .c_in(comb[30][17]), .S(S_s5_473), .c_out(C_s5_473));
FA FA_s5_480(.A(S_s6_482), .B(S_s6_481), .c_in(S_s6_480), .S(S_s5_480), .c_out(C_s5_480));
FA FA_s5_481(.A(C_s6_473), .B(C_s6_472), .c_in(C_s6_471), .S(S_s5_481), .c_out(C_s5_481));
FA FA_s5_482(.A(C_s6_470), .B(comb[26][22]), .c_in(comb[27][21]), .S(S_s5_482), .c_out(C_s5_482));
FA FA_s5_483(.A(comb[28][20]), .B(comb[29][19]), .c_in(comb[30][18]), .S(S_s5_483), .c_out(C_s5_483));
FA FA_s5_490(.A(S_s6_491), .B(S_s6_490), .c_in(C_s6_482), .S(S_s5_490), .c_out(C_s5_490));
FA FA_s5_491(.A(C_s6_481), .B(C_s6_480), .c_in(comb[24][25]), .S(S_s5_491), .c_out(C_s5_491));
FA FA_s5_492(.A(comb[25][24]), .B(comb[26][23]), .c_in(comb[27][22]), .S(S_s5_492), .c_out(C_s5_492));
FA FA_s5_493(.A(comb[28][21]), .B(comb[29][20]), .c_in(comb[30][19]), .S(S_s5_493), .c_out(C_s5_493));
FA FA_s5_500(.A(S_s6_500), .B(C_s6_491), .c_in(C_s6_490), .S(S_s5_500), .c_out(C_s5_500));
FA FA_s5_501(.A(comb[22][28]), .B(comb[23][27]), .c_in(comb[24][26]), .S(S_s5_501), .c_out(C_s5_501));
FA FA_s5_502(.A(comb[25][25]), .B(comb[26][24]), .c_in(comb[27][23]), .S(S_s5_502), .c_out(C_s5_502));
FA FA_s5_503(.A(comb[28][22]), .B(comb[29][21]), .c_in(comb[30][20]), .S(S_s5_503), .c_out(C_s5_503));
FA FA_s5_510(.A(C_s6_500), .B(comb[20][31]), .c_in(comb[21][30]), .S(S_s5_510), .c_out(C_s5_510));
FA FA_s5_511(.A(comb[22][29]), .B(comb[23][28]), .c_in(comb[24][27]), .S(S_s5_511), .c_out(C_s5_511));
FA FA_s5_512(.A(comb[25][26]), .B(comb[26][25]), .c_in(comb[27][24]), .S(S_s5_512), .c_out(C_s5_512));
FA FA_s5_513(.A(comb[28][23]), .B(comb[29][22]), .c_in(comb[30][21]), .S(S_s5_513), .c_out(C_s5_513));
FA FA_s5_520(.A(comb[21][31]), .B(comb[22][30]), .c_in(comb[23][29]), .S(S_s5_520), .c_out(C_s5_520));
FA FA_s5_521(.A(comb[24][28]), .B(comb[25][27]), .c_in(comb[26][26]), .S(S_s5_521), .c_out(C_s5_521));
FA FA_s5_522(.A(comb[27][25]), .B(comb[28][24]), .c_in(comb[29][23]), .S(S_s5_522), .c_out(C_s5_522));
FA FA_s5_530(.A(comb[22][31]), .B(comb[23][30]), .c_in(comb[24][29]), .S(S_s5_530), .c_out(C_s5_530));
FA FA_s5_531(.A(comb[25][28]), .B(comb[26][27]), .c_in(comb[27][26]), .S(S_s5_531), .c_out(C_s5_531));
FA FA_s5_540(.A(comb[23][31]), .B(comb[24][30]), .c_in(comb[25][29]), .S(S_s5_540), .c_out(C_s5_540));
// stage 5 end ======================================================================= 

// stage 4 begin ======================================================================= 
HA HA_s4_60(.A(comb[0][6]), .B(comb[1][5]), .S(S_s4_60), .c_out(C_s4_60));
FA FA_s4_70(.A(comb[0][7]), .B(comb[1][6]), .c_in(comb[2][5]), .S(S_s4_70), .c_out(C_s4_70));
HA HA_s4_71(.A(comb[3][4]), .B(comb[4][3]), .S(S_s4_71), .c_out(C_s4_71));
FA FA_s4_80(.A(comb[0][8]), .B(comb[1][7]), .c_in(comb[2][6]), .S(S_s4_80), .c_out(C_s4_80));
FA FA_s4_81(.A(comb[3][5]), .B(comb[4][4]), .c_in(comb[5][3]), .S(S_s4_81), .c_out(C_s4_81));
HA HA_s4_82(.A(comb[6][2]), .B(comb[7][1]), .S(S_s4_82), .c_out(C_s4_82));
FA FA_s4_90(.A(S_s5_90), .B(comb[2][7]), .c_in(comb[3][6]), .S(S_s4_90), .c_out(C_s4_90));
FA FA_s4_91(.A(comb[4][5]), .B(comb[5][4]), .c_in(comb[6][3]), .S(S_s4_91), .c_out(C_s4_91));
FA FA_s4_92(.A(comb[7][2]), .B(comb[8][1]), .c_in(comb[9][0]), .S(S_s4_92), .c_out(C_s4_92));
FA FA_s4_100(.A(S_s5_101), .B(S_s5_100), .c_in(C_s5_90), .S(S_s4_100), .c_out(C_s4_100));
FA FA_s4_101(.A(comb[5][5]), .B(comb[6][4]), .c_in(comb[7][3]), .S(S_s4_101), .c_out(C_s4_101));
FA FA_s4_102(.A(comb[8][2]), .B(comb[9][1]), .c_in(comb[10][0]), .S(S_s4_102), .c_out(C_s4_102));
FA FA_s4_110(.A(S_s5_112), .B(S_s5_111), .c_in(S_s5_110), .S(S_s4_110), .c_out(C_s4_110));
FA FA_s4_111(.A(C_s5_101), .B(C_s5_100), .c_in(comb[8][3]), .S(S_s4_111), .c_out(C_s4_111));
FA FA_s4_112(.A(comb[9][2]), .B(comb[10][1]), .c_in(comb[11][0]), .S(S_s4_112), .c_out(C_s4_112));
FA FA_s4_120(.A(S_s5_123), .B(S_s5_122), .c_in(S_s5_121), .S(S_s4_120), .c_out(C_s4_120));
FA FA_s4_121(.A(S_s5_120), .B(C_s5_112), .c_in(C_s5_111), .S(S_s4_121), .c_out(C_s4_121));
FA FA_s4_122(.A(C_s5_110), .B(comb[11][1]), .c_in(comb[12][0]), .S(S_s4_122), .c_out(C_s4_122));
FA FA_s4_130(.A(S_s5_133), .B(S_s5_132), .c_in(S_s5_131), .S(S_s4_130), .c_out(C_s4_130));
FA FA_s4_131(.A(S_s5_130), .B(C_s5_123), .c_in(C_s5_122), .S(S_s4_131), .c_out(C_s4_131));
FA FA_s4_132(.A(C_s5_121), .B(C_s5_120), .c_in(comb[13][0]), .S(S_s4_132), .c_out(C_s4_132));
FA FA_s4_140(.A(S_s5_143), .B(S_s5_142), .c_in(S_s5_141), .S(S_s4_140), .c_out(C_s4_140));
FA FA_s4_141(.A(S_s5_140), .B(C_s5_133), .c_in(C_s5_132), .S(S_s4_141), .c_out(C_s4_141));
FA FA_s4_142(.A(C_s5_131), .B(C_s5_130), .c_in(comb[14][0]), .S(S_s4_142), .c_out(C_s4_142));
FA FA_s4_150(.A(S_s5_153), .B(S_s5_152), .c_in(S_s5_151), .S(S_s4_150), .c_out(C_s4_150));
FA FA_s4_151(.A(S_s5_150), .B(C_s5_143), .c_in(C_s5_142), .S(S_s4_151), .c_out(C_s4_151));
FA FA_s4_152(.A(C_s5_141), .B(C_s5_140), .c_in(comb[15][0]), .S(S_s4_152), .c_out(C_s4_152));
FA FA_s4_160(.A(S_s5_163), .B(S_s5_162), .c_in(S_s5_161), .S(S_s4_160), .c_out(C_s4_160));
FA FA_s4_161(.A(S_s5_160), .B(C_s5_153), .c_in(C_s5_152), .S(S_s4_161), .c_out(C_s4_161));
FA FA_s4_162(.A(C_s5_151), .B(C_s5_150), .c_in(comb[16][0]), .S(S_s4_162), .c_out(C_s4_162));
FA FA_s4_170(.A(S_s5_173), .B(S_s5_172), .c_in(S_s5_171), .S(S_s4_170), .c_out(C_s4_170));
FA FA_s4_171(.A(S_s5_170), .B(C_s5_163), .c_in(C_s5_162), .S(S_s4_171), .c_out(C_s4_171));
FA FA_s4_172(.A(C_s5_161), .B(C_s5_160), .c_in(comb[17][0]), .S(S_s4_172), .c_out(C_s4_172));
FA FA_s4_180(.A(S_s5_183), .B(S_s5_182), .c_in(S_s5_181), .S(S_s4_180), .c_out(C_s4_180));
FA FA_s4_181(.A(S_s5_180), .B(C_s5_173), .c_in(C_s5_172), .S(S_s4_181), .c_out(C_s4_181));
FA FA_s4_182(.A(C_s5_171), .B(C_s5_170), .c_in(comb[18][0]), .S(S_s4_182), .c_out(C_s4_182));
FA FA_s4_190(.A(S_s5_193), .B(S_s5_192), .c_in(S_s5_191), .S(S_s4_190), .c_out(C_s4_190));
FA FA_s4_191(.A(S_s5_190), .B(C_s5_183), .c_in(C_s5_182), .S(S_s4_191), .c_out(C_s4_191));
FA FA_s4_192(.A(C_s5_181), .B(C_s5_180), .c_in(comb[19][0]), .S(S_s4_192), .c_out(C_s4_192));
FA FA_s4_200(.A(S_s5_203), .B(S_s5_202), .c_in(S_s5_201), .S(S_s4_200), .c_out(C_s4_200));
FA FA_s4_201(.A(S_s5_200), .B(C_s5_193), .c_in(C_s5_192), .S(S_s4_201), .c_out(C_s4_201));
FA FA_s4_202(.A(C_s5_191), .B(C_s5_190), .c_in(comb[20][0]), .S(S_s4_202), .c_out(C_s4_202));
FA FA_s4_210(.A(S_s5_213), .B(S_s5_212), .c_in(S_s5_211), .S(S_s4_210), .c_out(C_s4_210));
FA FA_s4_211(.A(S_s5_210), .B(C_s5_203), .c_in(C_s5_202), .S(S_s4_211), .c_out(C_s4_211));
FA FA_s4_212(.A(C_s5_201), .B(C_s5_200), .c_in(comb[21][0]), .S(S_s4_212), .c_out(C_s4_212));
FA FA_s4_220(.A(S_s5_223), .B(S_s5_222), .c_in(S_s5_221), .S(S_s4_220), .c_out(C_s4_220));
FA FA_s4_221(.A(S_s5_220), .B(C_s5_213), .c_in(C_s5_212), .S(S_s4_221), .c_out(C_s4_221));
FA FA_s4_222(.A(C_s5_211), .B(C_s5_210), .c_in(comb[22][0]), .S(S_s4_222), .c_out(C_s4_222));
FA FA_s4_230(.A(S_s5_233), .B(S_s5_232), .c_in(S_s5_231), .S(S_s4_230), .c_out(C_s4_230));
FA FA_s4_231(.A(S_s5_230), .B(C_s5_223), .c_in(C_s5_222), .S(S_s4_231), .c_out(C_s4_231));
FA FA_s4_232(.A(C_s5_221), .B(C_s5_220), .c_in(comb[23][0]), .S(S_s4_232), .c_out(C_s4_232));
FA FA_s4_240(.A(S_s5_243), .B(S_s5_242), .c_in(S_s5_241), .S(S_s4_240), .c_out(C_s4_240));
FA FA_s4_241(.A(S_s5_240), .B(C_s5_233), .c_in(C_s5_232), .S(S_s4_241), .c_out(C_s4_241));
FA FA_s4_242(.A(C_s5_231), .B(C_s5_230), .c_in(comb[24][0]), .S(S_s4_242), .c_out(C_s4_242));
FA FA_s4_250(.A(S_s5_253), .B(S_s5_252), .c_in(S_s5_251), .S(S_s4_250), .c_out(C_s4_250));
FA FA_s4_251(.A(S_s5_250), .B(C_s5_243), .c_in(C_s5_242), .S(S_s4_251), .c_out(C_s4_251));
FA FA_s4_252(.A(C_s5_241), .B(C_s5_240), .c_in(comb[25][0]), .S(S_s4_252), .c_out(C_s4_252));
FA FA_s4_260(.A(S_s5_263), .B(S_s5_262), .c_in(S_s5_261), .S(S_s4_260), .c_out(C_s4_260));
FA FA_s4_261(.A(S_s5_260), .B(C_s5_253), .c_in(C_s5_252), .S(S_s4_261), .c_out(C_s4_261));
FA FA_s4_262(.A(C_s5_251), .B(C_s5_250), .c_in(comb[26][0]), .S(S_s4_262), .c_out(C_s4_262));
FA FA_s4_270(.A(S_s5_273), .B(S_s5_272), .c_in(S_s5_271), .S(S_s4_270), .c_out(C_s4_270));
FA FA_s4_271(.A(S_s5_270), .B(C_s5_263), .c_in(C_s5_262), .S(S_s4_271), .c_out(C_s4_271));
FA FA_s4_272(.A(C_s5_261), .B(C_s5_260), .c_in(comb[27][0]), .S(S_s4_272), .c_out(C_s4_272));
FA FA_s4_280(.A(S_s5_283), .B(S_s5_282), .c_in(S_s5_281), .S(S_s4_280), .c_out(C_s4_280));
FA FA_s4_281(.A(S_s5_280), .B(C_s5_273), .c_in(C_s5_272), .S(S_s4_281), .c_out(C_s4_281));
FA FA_s4_282(.A(C_s5_271), .B(C_s5_270), .c_in(comb[28][0]), .S(S_s4_282), .c_out(C_s4_282));
FA FA_s4_290(.A(S_s5_293), .B(S_s5_292), .c_in(S_s5_291), .S(S_s4_290), .c_out(C_s4_290));
FA FA_s4_291(.A(S_s5_290), .B(C_s5_283), .c_in(C_s5_282), .S(S_s4_291), .c_out(C_s4_291));
FA FA_s4_292(.A(C_s5_281), .B(C_s5_280), .c_in(comb[29][0]), .S(S_s4_292), .c_out(C_s4_292));
FA FA_s4_300(.A(S_s5_303), .B(S_s5_302), .c_in(S_s5_301), .S(S_s4_300), .c_out(C_s4_300));
FA FA_s4_301(.A(S_s5_300), .B(C_s5_293), .c_in(C_s5_292), .S(S_s4_301), .c_out(C_s4_301));
FA FA_s4_302(.A(C_s5_291), .B(C_s5_290), .c_in(comb[30][0]), .S(S_s4_302), .c_out(C_s4_302));
FA FA_s4_310(.A(S_s5_313), .B(S_s5_312), .c_in(S_s5_311), .S(S_s4_310), .c_out(C_s4_310));
FA FA_s4_311(.A(S_s5_310), .B(C_s5_303), .c_in(C_s5_302), .S(S_s4_311), .c_out(C_s4_311));
FA FA_s4_312(.A(C_s5_301), .B(C_s5_300), .c_in(comb[31][0]), .S(S_s4_312), .c_out(C_s4_312));
FA FA_s4_320(.A(S_s5_323), .B(S_s5_322), .c_in(S_s5_321), .S(S_s4_320), .c_out(C_s4_320));
FA FA_s4_321(.A(S_s5_320), .B(C_s5_313), .c_in(C_s5_312), .S(S_s4_321), .c_out(C_s4_321));
FA FA_s4_322(.A(C_s5_311), .B(C_s5_310), .c_in(comb[31][1]), .S(S_s4_322), .c_out(C_s4_322));
FA FA_s4_330(.A(S_s5_333), .B(S_s5_332), .c_in(S_s5_331), .S(S_s4_330), .c_out(C_s4_330));
FA FA_s4_331(.A(S_s5_330), .B(C_s5_323), .c_in(C_s5_322), .S(S_s4_331), .c_out(C_s4_331));
FA FA_s4_332(.A(C_s5_321), .B(C_s5_320), .c_in(comb[31][2]), .S(S_s4_332), .c_out(C_s4_332));
FA FA_s4_340(.A(S_s5_343), .B(S_s5_342), .c_in(S_s5_341), .S(S_s4_340), .c_out(C_s4_340));
FA FA_s4_341(.A(S_s5_340), .B(C_s5_333), .c_in(C_s5_332), .S(S_s4_341), .c_out(C_s4_341));
FA FA_s4_342(.A(C_s5_331), .B(C_s5_330), .c_in(comb[31][3]), .S(S_s4_342), .c_out(C_s4_342));
FA FA_s4_350(.A(S_s5_353), .B(S_s5_352), .c_in(S_s5_351), .S(S_s4_350), .c_out(C_s4_350));
FA FA_s4_351(.A(S_s5_350), .B(C_s5_343), .c_in(C_s5_342), .S(S_s4_351), .c_out(C_s4_351));
FA FA_s4_352(.A(C_s5_341), .B(C_s5_340), .c_in(comb[31][4]), .S(S_s4_352), .c_out(C_s4_352));
FA FA_s4_360(.A(S_s5_363), .B(S_s5_362), .c_in(S_s5_361), .S(S_s4_360), .c_out(C_s4_360));
FA FA_s4_361(.A(S_s5_360), .B(C_s5_353), .c_in(C_s5_352), .S(S_s4_361), .c_out(C_s4_361));
FA FA_s4_362(.A(C_s5_351), .B(C_s5_350), .c_in(comb[31][5]), .S(S_s4_362), .c_out(C_s4_362));
FA FA_s4_370(.A(S_s5_373), .B(S_s5_372), .c_in(S_s5_371), .S(S_s4_370), .c_out(C_s4_370));
FA FA_s4_371(.A(S_s5_370), .B(C_s5_363), .c_in(C_s5_362), .S(S_s4_371), .c_out(C_s4_371));
FA FA_s4_372(.A(C_s5_361), .B(C_s5_360), .c_in(comb[31][6]), .S(S_s4_372), .c_out(C_s4_372));
FA FA_s4_380(.A(S_s5_383), .B(S_s5_382), .c_in(S_s5_381), .S(S_s4_380), .c_out(C_s4_380));
FA FA_s4_381(.A(S_s5_380), .B(C_s5_373), .c_in(C_s5_372), .S(S_s4_381), .c_out(C_s4_381));
FA FA_s4_382(.A(C_s5_371), .B(C_s5_370), .c_in(comb[31][7]), .S(S_s4_382), .c_out(C_s4_382));
FA FA_s4_390(.A(S_s5_393), .B(S_s5_392), .c_in(S_s5_391), .S(S_s4_390), .c_out(C_s4_390));
FA FA_s4_391(.A(S_s5_390), .B(C_s5_383), .c_in(C_s5_382), .S(S_s4_391), .c_out(C_s4_391));
FA FA_s4_392(.A(C_s5_381), .B(C_s5_380), .c_in(comb[31][8]), .S(S_s4_392), .c_out(C_s4_392));
FA FA_s4_400(.A(S_s5_403), .B(S_s5_402), .c_in(S_s5_401), .S(S_s4_400), .c_out(C_s4_400));
FA FA_s4_401(.A(S_s5_400), .B(C_s5_393), .c_in(C_s5_392), .S(S_s4_401), .c_out(C_s4_401));
FA FA_s4_402(.A(C_s5_391), .B(C_s5_390), .c_in(comb[31][9]), .S(S_s4_402), .c_out(C_s4_402));
FA FA_s4_410(.A(S_s5_413), .B(S_s5_412), .c_in(S_s5_411), .S(S_s4_410), .c_out(C_s4_410));
FA FA_s4_411(.A(S_s5_410), .B(C_s5_403), .c_in(C_s5_402), .S(S_s4_411), .c_out(C_s4_411));
FA FA_s4_412(.A(C_s5_401), .B(C_s5_400), .c_in(comb[31][10]), .S(S_s4_412), .c_out(C_s4_412));
FA FA_s4_420(.A(S_s5_423), .B(S_s5_422), .c_in(S_s5_421), .S(S_s4_420), .c_out(C_s4_420));
FA FA_s4_421(.A(S_s5_420), .B(C_s5_413), .c_in(C_s5_412), .S(S_s4_421), .c_out(C_s4_421));
FA FA_s4_422(.A(C_s5_411), .B(C_s5_410), .c_in(comb[31][11]), .S(S_s4_422), .c_out(C_s4_422));
FA FA_s4_430(.A(S_s5_433), .B(S_s5_432), .c_in(S_s5_431), .S(S_s4_430), .c_out(C_s4_430));
FA FA_s4_431(.A(S_s5_430), .B(C_s5_423), .c_in(C_s5_422), .S(S_s4_431), .c_out(C_s4_431));
FA FA_s4_432(.A(C_s5_421), .B(C_s5_420), .c_in(comb[31][12]), .S(S_s4_432), .c_out(C_s4_432));
FA FA_s4_440(.A(S_s5_443), .B(S_s5_442), .c_in(S_s5_441), .S(S_s4_440), .c_out(C_s4_440));
FA FA_s4_441(.A(S_s5_440), .B(C_s5_433), .c_in(C_s5_432), .S(S_s4_441), .c_out(C_s4_441));
FA FA_s4_442(.A(C_s5_431), .B(C_s5_430), .c_in(comb[31][13]), .S(S_s4_442), .c_out(C_s4_442));
FA FA_s4_450(.A(S_s5_453), .B(S_s5_452), .c_in(S_s5_451), .S(S_s4_450), .c_out(C_s4_450));
FA FA_s4_451(.A(S_s5_450), .B(C_s5_443), .c_in(C_s5_442), .S(S_s4_451), .c_out(C_s4_451));
FA FA_s4_452(.A(C_s5_441), .B(C_s5_440), .c_in(comb[31][14]), .S(S_s4_452), .c_out(C_s4_452));
FA FA_s4_460(.A(S_s5_463), .B(S_s5_462), .c_in(S_s5_461), .S(S_s4_460), .c_out(C_s4_460));
FA FA_s4_461(.A(S_s5_460), .B(C_s5_453), .c_in(C_s5_452), .S(S_s4_461), .c_out(C_s4_461));
FA FA_s4_462(.A(C_s5_451), .B(C_s5_450), .c_in(comb[31][15]), .S(S_s4_462), .c_out(C_s4_462));
FA FA_s4_470(.A(S_s5_473), .B(S_s5_472), .c_in(S_s5_471), .S(S_s4_470), .c_out(C_s4_470));
FA FA_s4_471(.A(S_s5_470), .B(C_s5_463), .c_in(C_s5_462), .S(S_s4_471), .c_out(C_s4_471));
FA FA_s4_472(.A(C_s5_461), .B(C_s5_460), .c_in(comb[31][16]), .S(S_s4_472), .c_out(C_s4_472));
FA FA_s4_480(.A(S_s5_483), .B(S_s5_482), .c_in(S_s5_481), .S(S_s4_480), .c_out(C_s4_480));
FA FA_s4_481(.A(S_s5_480), .B(C_s5_473), .c_in(C_s5_472), .S(S_s4_481), .c_out(C_s4_481));
FA FA_s4_482(.A(C_s5_471), .B(C_s5_470), .c_in(comb[31][17]), .S(S_s4_482), .c_out(C_s4_482));
FA FA_s4_490(.A(S_s5_493), .B(S_s5_492), .c_in(S_s5_491), .S(S_s4_490), .c_out(C_s4_490));
FA FA_s4_491(.A(S_s5_490), .B(C_s5_483), .c_in(C_s5_482), .S(S_s4_491), .c_out(C_s4_491));
FA FA_s4_492(.A(C_s5_481), .B(C_s5_480), .c_in(comb[31][18]), .S(S_s4_492), .c_out(C_s4_492));
FA FA_s4_500(.A(S_s5_503), .B(S_s5_502), .c_in(S_s5_501), .S(S_s4_500), .c_out(C_s4_500));
FA FA_s4_501(.A(S_s5_500), .B(C_s5_493), .c_in(C_s5_492), .S(S_s4_501), .c_out(C_s4_501));
FA FA_s4_502(.A(C_s5_491), .B(C_s5_490), .c_in(comb[31][19]), .S(S_s4_502), .c_out(C_s4_502));
FA FA_s4_510(.A(S_s5_513), .B(S_s5_512), .c_in(S_s5_511), .S(S_s4_510), .c_out(C_s4_510));
FA FA_s4_511(.A(S_s5_510), .B(C_s5_503), .c_in(C_s5_502), .S(S_s4_511), .c_out(C_s4_511));
FA FA_s4_512(.A(C_s5_501), .B(C_s5_500), .c_in(comb[31][20]), .S(S_s4_512), .c_out(C_s4_512));
FA FA_s4_520(.A(S_s5_522), .B(S_s5_521), .c_in(S_s5_520), .S(S_s4_520), .c_out(C_s4_520));
FA FA_s4_521(.A(C_s5_513), .B(C_s5_512), .c_in(C_s5_511), .S(S_s4_521), .c_out(C_s4_521));
FA FA_s4_522(.A(C_s5_510), .B(comb[30][22]), .c_in(comb[31][21]), .S(S_s4_522), .c_out(C_s4_522));
FA FA_s4_530(.A(S_s5_531), .B(S_s5_530), .c_in(C_s5_522), .S(S_s4_530), .c_out(C_s4_530));
FA FA_s4_531(.A(C_s5_521), .B(C_s5_520), .c_in(comb[28][25]), .S(S_s4_531), .c_out(C_s4_531));
FA FA_s4_532(.A(comb[29][24]), .B(comb[30][23]), .c_in(comb[31][22]), .S(S_s4_532), .c_out(C_s4_532));
FA FA_s4_540(.A(S_s5_540), .B(C_s5_531), .c_in(C_s5_530), .S(S_s4_540), .c_out(C_s4_540));
FA FA_s4_541(.A(comb[26][28]), .B(comb[27][27]), .c_in(comb[28][26]), .S(S_s4_541), .c_out(C_s4_541));
FA FA_s4_542(.A(comb[29][25]), .B(comb[30][24]), .c_in(comb[31][23]), .S(S_s4_542), .c_out(C_s4_542));
FA FA_s4_550(.A(C_s5_540), .B(comb[24][31]), .c_in(comb[25][30]), .S(S_s4_550), .c_out(C_s4_550));
FA FA_s4_551(.A(comb[26][29]), .B(comb[27][28]), .c_in(comb[28][27]), .S(S_s4_551), .c_out(C_s4_551));
FA FA_s4_552(.A(comb[29][26]), .B(comb[30][25]), .c_in(comb[31][24]), .S(S_s4_552), .c_out(C_s4_552));
FA FA_s4_560(.A(comb[25][31]), .B(comb[26][30]), .c_in(comb[27][29]), .S(S_s4_560), .c_out(C_s4_560));
FA FA_s4_561(.A(comb[28][28]), .B(comb[29][27]), .c_in(comb[30][26]), .S(S_s4_561), .c_out(C_s4_561));
FA FA_s4_570(.A(comb[26][31]), .B(comb[27][30]), .c_in(comb[28][29]), .S(S_s4_570), .c_out(C_s4_570));
// stage 4 end ======================================================================= 

// stage 3 begin ======================================================================= 
HA HA_s3_40(.A(comb[0][4]), .B(comb[1][3]), .S(S_s3_40), .c_out(C_s3_40));
FA FA_s3_50(.A(comb[0][5]), .B(comb[1][4]), .c_in(comb[2][3]), .S(S_s3_50), .c_out(C_s3_50));
HA HA_s3_51(.A(comb[3][2]), .B(comb[4][1]), .S(S_s3_51), .c_out(C_s3_51));
FA FA_s3_60(.A(S_s4_60), .B(comb[2][4]), .c_in(comb[3][3]), .S(S_s3_60), .c_out(C_s3_60));
FA FA_s3_61(.A(comb[4][2]), .B(comb[5][1]), .c_in(comb[6][0]), .S(S_s3_61), .c_out(C_s3_61));
FA FA_s3_70(.A(S_s4_71), .B(S_s4_70), .c_in(C_s4_60), .S(S_s3_70), .c_out(C_s3_70));
FA FA_s3_71(.A(comb[5][2]), .B(comb[6][1]), .c_in(comb[7][0]), .S(S_s3_71), .c_out(C_s3_71));
FA FA_s3_80(.A(S_s4_82), .B(S_s4_81), .c_in(S_s4_80), .S(S_s3_80), .c_out(C_s3_80));
FA FA_s3_81(.A(C_s4_71), .B(C_s4_70), .c_in(comb[8][0]), .S(S_s3_81), .c_out(C_s3_81));
FA FA_s3_90(.A(S_s4_92), .B(S_s4_91), .c_in(S_s4_90), .S(S_s3_90), .c_out(C_s3_90));
FA FA_s3_91(.A(C_s4_82), .B(C_s4_81), .c_in(C_s4_80), .S(S_s3_91), .c_out(C_s3_91));
FA FA_s3_100(.A(S_s4_102), .B(S_s4_101), .c_in(S_s4_100), .S(S_s3_100), .c_out(C_s3_100));
FA FA_s3_101(.A(C_s4_92), .B(C_s4_91), .c_in(C_s4_90), .S(S_s3_101), .c_out(C_s3_101));
FA FA_s3_110(.A(S_s4_112), .B(S_s4_111), .c_in(S_s4_110), .S(S_s3_110), .c_out(C_s3_110));
FA FA_s3_111(.A(C_s4_102), .B(C_s4_101), .c_in(C_s4_100), .S(S_s3_111), .c_out(C_s3_111));
FA FA_s3_120(.A(S_s4_122), .B(S_s4_121), .c_in(S_s4_120), .S(S_s3_120), .c_out(C_s3_120));
FA FA_s3_121(.A(C_s4_112), .B(C_s4_111), .c_in(C_s4_110), .S(S_s3_121), .c_out(C_s3_121));
FA FA_s3_130(.A(S_s4_132), .B(S_s4_131), .c_in(S_s4_130), .S(S_s3_130), .c_out(C_s3_130));
FA FA_s3_131(.A(C_s4_122), .B(C_s4_121), .c_in(C_s4_120), .S(S_s3_131), .c_out(C_s3_131));
FA FA_s3_140(.A(S_s4_142), .B(S_s4_141), .c_in(S_s4_140), .S(S_s3_140), .c_out(C_s3_140));
FA FA_s3_141(.A(C_s4_132), .B(C_s4_131), .c_in(C_s4_130), .S(S_s3_141), .c_out(C_s3_141));
FA FA_s3_150(.A(S_s4_152), .B(S_s4_151), .c_in(S_s4_150), .S(S_s3_150), .c_out(C_s3_150));
FA FA_s3_151(.A(C_s4_142), .B(C_s4_141), .c_in(C_s4_140), .S(S_s3_151), .c_out(C_s3_151));
FA FA_s3_160(.A(S_s4_162), .B(S_s4_161), .c_in(S_s4_160), .S(S_s3_160), .c_out(C_s3_160));
FA FA_s3_161(.A(C_s4_152), .B(C_s4_151), .c_in(C_s4_150), .S(S_s3_161), .c_out(C_s3_161));
FA FA_s3_170(.A(S_s4_172), .B(S_s4_171), .c_in(S_s4_170), .S(S_s3_170), .c_out(C_s3_170));
FA FA_s3_171(.A(C_s4_162), .B(C_s4_161), .c_in(C_s4_160), .S(S_s3_171), .c_out(C_s3_171));
FA FA_s3_180(.A(S_s4_182), .B(S_s4_181), .c_in(S_s4_180), .S(S_s3_180), .c_out(C_s3_180));
FA FA_s3_181(.A(C_s4_172), .B(C_s4_171), .c_in(C_s4_170), .S(S_s3_181), .c_out(C_s3_181));
FA FA_s3_190(.A(S_s4_192), .B(S_s4_191), .c_in(S_s4_190), .S(S_s3_190), .c_out(C_s3_190));
FA FA_s3_191(.A(C_s4_182), .B(C_s4_181), .c_in(C_s4_180), .S(S_s3_191), .c_out(C_s3_191));
FA FA_s3_200(.A(S_s4_202), .B(S_s4_201), .c_in(S_s4_200), .S(S_s3_200), .c_out(C_s3_200));
FA FA_s3_201(.A(C_s4_192), .B(C_s4_191), .c_in(C_s4_190), .S(S_s3_201), .c_out(C_s3_201));
FA FA_s3_210(.A(S_s4_212), .B(S_s4_211), .c_in(S_s4_210), .S(S_s3_210), .c_out(C_s3_210));
FA FA_s3_211(.A(C_s4_202), .B(C_s4_201), .c_in(C_s4_200), .S(S_s3_211), .c_out(C_s3_211));
FA FA_s3_220(.A(S_s4_222), .B(S_s4_221), .c_in(S_s4_220), .S(S_s3_220), .c_out(C_s3_220));
FA FA_s3_221(.A(C_s4_212), .B(C_s4_211), .c_in(C_s4_210), .S(S_s3_221), .c_out(C_s3_221));
FA FA_s3_230(.A(S_s4_232), .B(S_s4_231), .c_in(S_s4_230), .S(S_s3_230), .c_out(C_s3_230));
FA FA_s3_231(.A(C_s4_222), .B(C_s4_221), .c_in(C_s4_220), .S(S_s3_231), .c_out(C_s3_231));
FA FA_s3_240(.A(S_s4_242), .B(S_s4_241), .c_in(S_s4_240), .S(S_s3_240), .c_out(C_s3_240));
FA FA_s3_241(.A(C_s4_232), .B(C_s4_231), .c_in(C_s4_230), .S(S_s3_241), .c_out(C_s3_241));
FA FA_s3_250(.A(S_s4_252), .B(S_s4_251), .c_in(S_s4_250), .S(S_s3_250), .c_out(C_s3_250));
FA FA_s3_251(.A(C_s4_242), .B(C_s4_241), .c_in(C_s4_240), .S(S_s3_251), .c_out(C_s3_251));
FA FA_s3_260(.A(S_s4_262), .B(S_s4_261), .c_in(S_s4_260), .S(S_s3_260), .c_out(C_s3_260));
FA FA_s3_261(.A(C_s4_252), .B(C_s4_251), .c_in(C_s4_250), .S(S_s3_261), .c_out(C_s3_261));
FA FA_s3_270(.A(S_s4_272), .B(S_s4_271), .c_in(S_s4_270), .S(S_s3_270), .c_out(C_s3_270));
FA FA_s3_271(.A(C_s4_262), .B(C_s4_261), .c_in(C_s4_260), .S(S_s3_271), .c_out(C_s3_271));
FA FA_s3_280(.A(S_s4_282), .B(S_s4_281), .c_in(S_s4_280), .S(S_s3_280), .c_out(C_s3_280));
FA FA_s3_281(.A(C_s4_272), .B(C_s4_271), .c_in(C_s4_270), .S(S_s3_281), .c_out(C_s3_281));
FA FA_s3_290(.A(S_s4_292), .B(S_s4_291), .c_in(S_s4_290), .S(S_s3_290), .c_out(C_s3_290));
FA FA_s3_291(.A(C_s4_282), .B(C_s4_281), .c_in(C_s4_280), .S(S_s3_291), .c_out(C_s3_291));
FA FA_s3_300(.A(S_s4_302), .B(S_s4_301), .c_in(S_s4_300), .S(S_s3_300), .c_out(C_s3_300));
FA FA_s3_301(.A(C_s4_292), .B(C_s4_291), .c_in(C_s4_290), .S(S_s3_301), .c_out(C_s3_301));
FA FA_s3_310(.A(S_s4_312), .B(S_s4_311), .c_in(S_s4_310), .S(S_s3_310), .c_out(C_s3_310));
FA FA_s3_311(.A(C_s4_302), .B(C_s4_301), .c_in(C_s4_300), .S(S_s3_311), .c_out(C_s3_311));
FA FA_s3_320(.A(S_s4_322), .B(S_s4_321), .c_in(S_s4_320), .S(S_s3_320), .c_out(C_s3_320));
FA FA_s3_321(.A(C_s4_312), .B(C_s4_311), .c_in(C_s4_310), .S(S_s3_321), .c_out(C_s3_321));
FA FA_s3_330(.A(S_s4_332), .B(S_s4_331), .c_in(S_s4_330), .S(S_s3_330), .c_out(C_s3_330));
FA FA_s3_331(.A(C_s4_322), .B(C_s4_321), .c_in(C_s4_320), .S(S_s3_331), .c_out(C_s3_331));
FA FA_s3_340(.A(S_s4_342), .B(S_s4_341), .c_in(S_s4_340), .S(S_s3_340), .c_out(C_s3_340));
FA FA_s3_341(.A(C_s4_332), .B(C_s4_331), .c_in(C_s4_330), .S(S_s3_341), .c_out(C_s3_341));
FA FA_s3_350(.A(S_s4_352), .B(S_s4_351), .c_in(S_s4_350), .S(S_s3_350), .c_out(C_s3_350));
FA FA_s3_351(.A(C_s4_342), .B(C_s4_341), .c_in(C_s4_340), .S(S_s3_351), .c_out(C_s3_351));
FA FA_s3_360(.A(S_s4_362), .B(S_s4_361), .c_in(S_s4_360), .S(S_s3_360), .c_out(C_s3_360));
FA FA_s3_361(.A(C_s4_352), .B(C_s4_351), .c_in(C_s4_350), .S(S_s3_361), .c_out(C_s3_361));
FA FA_s3_370(.A(S_s4_372), .B(S_s4_371), .c_in(S_s4_370), .S(S_s3_370), .c_out(C_s3_370));
FA FA_s3_371(.A(C_s4_362), .B(C_s4_361), .c_in(C_s4_360), .S(S_s3_371), .c_out(C_s3_371));
FA FA_s3_380(.A(S_s4_382), .B(S_s4_381), .c_in(S_s4_380), .S(S_s3_380), .c_out(C_s3_380));
FA FA_s3_381(.A(C_s4_372), .B(C_s4_371), .c_in(C_s4_370), .S(S_s3_381), .c_out(C_s3_381));
FA FA_s3_390(.A(S_s4_392), .B(S_s4_391), .c_in(S_s4_390), .S(S_s3_390), .c_out(C_s3_390));
FA FA_s3_391(.A(C_s4_382), .B(C_s4_381), .c_in(C_s4_380), .S(S_s3_391), .c_out(C_s3_391));
FA FA_s3_400(.A(S_s4_402), .B(S_s4_401), .c_in(S_s4_400), .S(S_s3_400), .c_out(C_s3_400));
FA FA_s3_401(.A(C_s4_392), .B(C_s4_391), .c_in(C_s4_390), .S(S_s3_401), .c_out(C_s3_401));
FA FA_s3_410(.A(S_s4_412), .B(S_s4_411), .c_in(S_s4_410), .S(S_s3_410), .c_out(C_s3_410));
FA FA_s3_411(.A(C_s4_402), .B(C_s4_401), .c_in(C_s4_400), .S(S_s3_411), .c_out(C_s3_411));
FA FA_s3_420(.A(S_s4_422), .B(S_s4_421), .c_in(S_s4_420), .S(S_s3_420), .c_out(C_s3_420));
FA FA_s3_421(.A(C_s4_412), .B(C_s4_411), .c_in(C_s4_410), .S(S_s3_421), .c_out(C_s3_421));
FA FA_s3_430(.A(S_s4_432), .B(S_s4_431), .c_in(S_s4_430), .S(S_s3_430), .c_out(C_s3_430));
FA FA_s3_431(.A(C_s4_422), .B(C_s4_421), .c_in(C_s4_420), .S(S_s3_431), .c_out(C_s3_431));
FA FA_s3_440(.A(S_s4_442), .B(S_s4_441), .c_in(S_s4_440), .S(S_s3_440), .c_out(C_s3_440));
FA FA_s3_441(.A(C_s4_432), .B(C_s4_431), .c_in(C_s4_430), .S(S_s3_441), .c_out(C_s3_441));
FA FA_s3_450(.A(S_s4_452), .B(S_s4_451), .c_in(S_s4_450), .S(S_s3_450), .c_out(C_s3_450));
FA FA_s3_451(.A(C_s4_442), .B(C_s4_441), .c_in(C_s4_440), .S(S_s3_451), .c_out(C_s3_451));
FA FA_s3_460(.A(S_s4_462), .B(S_s4_461), .c_in(S_s4_460), .S(S_s3_460), .c_out(C_s3_460));
FA FA_s3_461(.A(C_s4_452), .B(C_s4_451), .c_in(C_s4_450), .S(S_s3_461), .c_out(C_s3_461));
FA FA_s3_470(.A(S_s4_472), .B(S_s4_471), .c_in(S_s4_470), .S(S_s3_470), .c_out(C_s3_470));
FA FA_s3_471(.A(C_s4_462), .B(C_s4_461), .c_in(C_s4_460), .S(S_s3_471), .c_out(C_s3_471));
FA FA_s3_480(.A(S_s4_482), .B(S_s4_481), .c_in(S_s4_480), .S(S_s3_480), .c_out(C_s3_480));
FA FA_s3_481(.A(C_s4_472), .B(C_s4_471), .c_in(C_s4_470), .S(S_s3_481), .c_out(C_s3_481));
FA FA_s3_490(.A(S_s4_492), .B(S_s4_491), .c_in(S_s4_490), .S(S_s3_490), .c_out(C_s3_490));
FA FA_s3_491(.A(C_s4_482), .B(C_s4_481), .c_in(C_s4_480), .S(S_s3_491), .c_out(C_s3_491));
FA FA_s3_500(.A(S_s4_502), .B(S_s4_501), .c_in(S_s4_500), .S(S_s3_500), .c_out(C_s3_500));
FA FA_s3_501(.A(C_s4_492), .B(C_s4_491), .c_in(C_s4_490), .S(S_s3_501), .c_out(C_s3_501));
FA FA_s3_510(.A(S_s4_512), .B(S_s4_511), .c_in(S_s4_510), .S(S_s3_510), .c_out(C_s3_510));
FA FA_s3_511(.A(C_s4_502), .B(C_s4_501), .c_in(C_s4_500), .S(S_s3_511), .c_out(C_s3_511));
FA FA_s3_520(.A(S_s4_522), .B(S_s4_521), .c_in(S_s4_520), .S(S_s3_520), .c_out(C_s3_520));
FA FA_s3_521(.A(C_s4_512), .B(C_s4_511), .c_in(C_s4_510), .S(S_s3_521), .c_out(C_s3_521));
FA FA_s3_530(.A(S_s4_532), .B(S_s4_531), .c_in(S_s4_530), .S(S_s3_530), .c_out(C_s3_530));
FA FA_s3_531(.A(C_s4_522), .B(C_s4_521), .c_in(C_s4_520), .S(S_s3_531), .c_out(C_s3_531));
FA FA_s3_540(.A(S_s4_542), .B(S_s4_541), .c_in(S_s4_540), .S(S_s3_540), .c_out(C_s3_540));
FA FA_s3_541(.A(C_s4_532), .B(C_s4_531), .c_in(C_s4_530), .S(S_s3_541), .c_out(C_s3_541));
FA FA_s3_550(.A(S_s4_552), .B(S_s4_551), .c_in(S_s4_550), .S(S_s3_550), .c_out(C_s3_550));
FA FA_s3_551(.A(C_s4_542), .B(C_s4_541), .c_in(C_s4_540), .S(S_s3_551), .c_out(C_s3_551));
FA FA_s3_560(.A(S_s4_561), .B(S_s4_560), .c_in(C_s4_552), .S(S_s3_560), .c_out(C_s3_560));
FA FA_s3_561(.A(C_s4_551), .B(C_s4_550), .c_in(comb[31][25]), .S(S_s3_561), .c_out(C_s3_561));
FA FA_s3_570(.A(S_s4_570), .B(C_s4_561), .c_in(C_s4_560), .S(S_s3_570), .c_out(C_s3_570));
FA FA_s3_571(.A(comb[29][28]), .B(comb[30][27]), .c_in(comb[31][26]), .S(S_s3_571), .c_out(C_s3_571));
FA FA_s3_580(.A(C_s4_570), .B(comb[27][31]), .c_in(comb[28][30]), .S(S_s3_580), .c_out(C_s3_580));
FA FA_s3_581(.A(comb[29][29]), .B(comb[30][28]), .c_in(comb[31][27]), .S(S_s3_581), .c_out(C_s3_581));
FA FA_s3_590(.A(comb[28][31]), .B(comb[29][30]), .c_in(comb[30][29]), .S(S_s3_590), .c_out(C_s3_590));
// stage 3 end ======================================================================= 

// stage 2 begin ======================================================================= 
HA HA_s2_30(.A(comb[0][3]), .B(comb[1][2]), .S(S_s2_30), .c_out(C_s2_30));
FA FA_s2_40(.A(S_s3_40), .B(comb[2][2]), .c_in(comb[3][1]), .S(S_s2_40), .c_out(C_s2_40));
FA FA_s2_50(.A(S_s3_51), .B(S_s3_50), .c_in(C_s3_40), .S(S_s2_50), .c_out(C_s2_50));
FA FA_s2_60(.A(S_s3_61), .B(S_s3_60), .c_in(C_s3_51), .S(S_s2_60), .c_out(C_s2_60));
FA FA_s2_70(.A(S_s3_71), .B(S_s3_70), .c_in(C_s3_61), .S(S_s2_70), .c_out(C_s2_70));
FA FA_s2_80(.A(S_s3_81), .B(S_s3_80), .c_in(C_s3_71), .S(S_s2_80), .c_out(C_s2_80));
FA FA_s2_90(.A(S_s3_91), .B(S_s3_90), .c_in(C_s3_81), .S(S_s2_90), .c_out(C_s2_90));
FA FA_s2_100(.A(S_s3_101), .B(S_s3_100), .c_in(C_s3_91), .S(S_s2_100), .c_out(C_s2_100));
FA FA_s2_110(.A(S_s3_111), .B(S_s3_110), .c_in(C_s3_101), .S(S_s2_110), .c_out(C_s2_110));
FA FA_s2_120(.A(S_s3_121), .B(S_s3_120), .c_in(C_s3_111), .S(S_s2_120), .c_out(C_s2_120));
FA FA_s2_130(.A(S_s3_131), .B(S_s3_130), .c_in(C_s3_121), .S(S_s2_130), .c_out(C_s2_130));
FA FA_s2_140(.A(S_s3_141), .B(S_s3_140), .c_in(C_s3_131), .S(S_s2_140), .c_out(C_s2_140));
FA FA_s2_150(.A(S_s3_151), .B(S_s3_150), .c_in(C_s3_141), .S(S_s2_150), .c_out(C_s2_150));
FA FA_s2_160(.A(S_s3_161), .B(S_s3_160), .c_in(C_s3_151), .S(S_s2_160), .c_out(C_s2_160));
FA FA_s2_170(.A(S_s3_171), .B(S_s3_170), .c_in(C_s3_161), .S(S_s2_170), .c_out(C_s2_170));
FA FA_s2_180(.A(S_s3_181), .B(S_s3_180), .c_in(C_s3_171), .S(S_s2_180), .c_out(C_s2_180));
FA FA_s2_190(.A(S_s3_191), .B(S_s3_190), .c_in(C_s3_181), .S(S_s2_190), .c_out(C_s2_190));
FA FA_s2_200(.A(S_s3_201), .B(S_s3_200), .c_in(C_s3_191), .S(S_s2_200), .c_out(C_s2_200));
FA FA_s2_210(.A(S_s3_211), .B(S_s3_210), .c_in(C_s3_201), .S(S_s2_210), .c_out(C_s2_210));
FA FA_s2_220(.A(S_s3_221), .B(S_s3_220), .c_in(C_s3_211), .S(S_s2_220), .c_out(C_s2_220));
FA FA_s2_230(.A(S_s3_231), .B(S_s3_230), .c_in(C_s3_221), .S(S_s2_230), .c_out(C_s2_230));
FA FA_s2_240(.A(S_s3_241), .B(S_s3_240), .c_in(C_s3_231), .S(S_s2_240), .c_out(C_s2_240));
FA FA_s2_250(.A(S_s3_251), .B(S_s3_250), .c_in(C_s3_241), .S(S_s2_250), .c_out(C_s2_250));
FA FA_s2_260(.A(S_s3_261), .B(S_s3_260), .c_in(C_s3_251), .S(S_s2_260), .c_out(C_s2_260));
FA FA_s2_270(.A(S_s3_271), .B(S_s3_270), .c_in(C_s3_261), .S(S_s2_270), .c_out(C_s2_270));
FA FA_s2_280(.A(S_s3_281), .B(S_s3_280), .c_in(C_s3_271), .S(S_s2_280), .c_out(C_s2_280));
FA FA_s2_290(.A(S_s3_291), .B(S_s3_290), .c_in(C_s3_281), .S(S_s2_290), .c_out(C_s2_290));
FA FA_s2_300(.A(S_s3_301), .B(S_s3_300), .c_in(C_s3_291), .S(S_s2_300), .c_out(C_s2_300));
FA FA_s2_310(.A(S_s3_311), .B(S_s3_310), .c_in(C_s3_301), .S(S_s2_310), .c_out(C_s2_310));
FA FA_s2_320(.A(S_s3_321), .B(S_s3_320), .c_in(C_s3_311), .S(S_s2_320), .c_out(C_s2_320));
FA FA_s2_330(.A(S_s3_331), .B(S_s3_330), .c_in(C_s3_321), .S(S_s2_330), .c_out(C_s2_330));
FA FA_s2_340(.A(S_s3_341), .B(S_s3_340), .c_in(C_s3_331), .S(S_s2_340), .c_out(C_s2_340));
FA FA_s2_350(.A(S_s3_351), .B(S_s3_350), .c_in(C_s3_341), .S(S_s2_350), .c_out(C_s2_350));
FA FA_s2_360(.A(S_s3_361), .B(S_s3_360), .c_in(C_s3_351), .S(S_s2_360), .c_out(C_s2_360));
FA FA_s2_370(.A(S_s3_371), .B(S_s3_370), .c_in(C_s3_361), .S(S_s2_370), .c_out(C_s2_370));
FA FA_s2_380(.A(S_s3_381), .B(S_s3_380), .c_in(C_s3_371), .S(S_s2_380), .c_out(C_s2_380));
FA FA_s2_390(.A(S_s3_391), .B(S_s3_390), .c_in(C_s3_381), .S(S_s2_390), .c_out(C_s2_390));
FA FA_s2_400(.A(S_s3_401), .B(S_s3_400), .c_in(C_s3_391), .S(S_s2_400), .c_out(C_s2_400));
FA FA_s2_410(.A(S_s3_411), .B(S_s3_410), .c_in(C_s3_401), .S(S_s2_410), .c_out(C_s2_410));
FA FA_s2_420(.A(S_s3_421), .B(S_s3_420), .c_in(C_s3_411), .S(S_s2_420), .c_out(C_s2_420));
FA FA_s2_430(.A(S_s3_431), .B(S_s3_430), .c_in(C_s3_421), .S(S_s2_430), .c_out(C_s2_430));
FA FA_s2_440(.A(S_s3_441), .B(S_s3_440), .c_in(C_s3_431), .S(S_s2_440), .c_out(C_s2_440));
FA FA_s2_450(.A(S_s3_451), .B(S_s3_450), .c_in(C_s3_441), .S(S_s2_450), .c_out(C_s2_450));
FA FA_s2_460(.A(S_s3_461), .B(S_s3_460), .c_in(C_s3_451), .S(S_s2_460), .c_out(C_s2_460));
FA FA_s2_470(.A(S_s3_471), .B(S_s3_470), .c_in(C_s3_461), .S(S_s2_470), .c_out(C_s2_470));
FA FA_s2_480(.A(S_s3_481), .B(S_s3_480), .c_in(C_s3_471), .S(S_s2_480), .c_out(C_s2_480));
FA FA_s2_490(.A(S_s3_491), .B(S_s3_490), .c_in(C_s3_481), .S(S_s2_490), .c_out(C_s2_490));
FA FA_s2_500(.A(S_s3_501), .B(S_s3_500), .c_in(C_s3_491), .S(S_s2_500), .c_out(C_s2_500));
FA FA_s2_510(.A(S_s3_511), .B(S_s3_510), .c_in(C_s3_501), .S(S_s2_510), .c_out(C_s2_510));
FA FA_s2_520(.A(S_s3_521), .B(S_s3_520), .c_in(C_s3_511), .S(S_s2_520), .c_out(C_s2_520));
FA FA_s2_530(.A(S_s3_531), .B(S_s3_530), .c_in(C_s3_521), .S(S_s2_530), .c_out(C_s2_530));
FA FA_s2_540(.A(S_s3_541), .B(S_s3_540), .c_in(C_s3_531), .S(S_s2_540), .c_out(C_s2_540));
FA FA_s2_550(.A(S_s3_551), .B(S_s3_550), .c_in(C_s3_541), .S(S_s2_550), .c_out(C_s2_550));
FA FA_s2_560(.A(S_s3_561), .B(S_s3_560), .c_in(C_s3_551), .S(S_s2_560), .c_out(C_s2_560));
FA FA_s2_570(.A(S_s3_571), .B(S_s3_570), .c_in(C_s3_561), .S(S_s2_570), .c_out(C_s2_570));
FA FA_s2_580(.A(S_s3_581), .B(S_s3_580), .c_in(C_s3_571), .S(S_s2_580), .c_out(C_s2_580));
FA FA_s2_590(.A(S_s3_590), .B(C_s3_581), .c_in(C_s3_580), .S(S_s2_590), .c_out(C_s2_590));
FA FA_s2_600(.A(C_s3_590), .B(comb[29][31]), .c_in(comb[30][30]), .S(S_s2_600), .c_out(C_s2_600));
// stage 2 end ======================================================================= 

// stage 1 begin ======================================================================= 
HA HA_s1_20(.A(comb[0][2]), .B(comb[1][1]), .S(S_s1_20), .c_out(C_s1_20));
FA FA_s1_30(.A(S_s2_30), .B(comb[2][1]), .c_in(comb[3][0]), .S(S_s1_30), .c_out(C_s1_30));
FA FA_s1_40(.A(S_s2_40), .B(C_s2_30), .c_in(comb[4][0]), .S(S_s1_40), .c_out(C_s1_40));
FA FA_s1_50(.A(S_s2_50), .B(C_s2_40), .c_in(comb[5][0]), .S(S_s1_50), .c_out(C_s1_50));
FA FA_s1_60(.A(S_s2_60), .B(C_s2_50), .c_in(C_s3_50), .S(S_s1_60), .c_out(C_s1_60));
FA FA_s1_70(.A(S_s2_70), .B(C_s2_60), .c_in(C_s3_60), .S(S_s1_70), .c_out(C_s1_70));
FA FA_s1_80(.A(S_s2_80), .B(C_s2_70), .c_in(C_s3_70), .S(S_s1_80), .c_out(C_s1_80));
FA FA_s1_90(.A(S_s2_90), .B(C_s2_80), .c_in(C_s3_80), .S(S_s1_90), .c_out(C_s1_90));
FA FA_s1_100(.A(S_s2_100), .B(C_s2_90), .c_in(C_s3_90), .S(S_s1_100), .c_out(C_s1_100));
FA FA_s1_110(.A(S_s2_110), .B(C_s2_100), .c_in(C_s3_100), .S(S_s1_110), .c_out(C_s1_110));
FA FA_s1_120(.A(S_s2_120), .B(C_s2_110), .c_in(C_s3_110), .S(S_s1_120), .c_out(C_s1_120));
FA FA_s1_130(.A(S_s2_130), .B(C_s2_120), .c_in(C_s3_120), .S(S_s1_130), .c_out(C_s1_130));
FA FA_s1_140(.A(S_s2_140), .B(C_s2_130), .c_in(C_s3_130), .S(S_s1_140), .c_out(C_s1_140));
FA FA_s1_150(.A(S_s2_150), .B(C_s2_140), .c_in(C_s3_140), .S(S_s1_150), .c_out(C_s1_150));
FA FA_s1_160(.A(S_s2_160), .B(C_s2_150), .c_in(C_s3_150), .S(S_s1_160), .c_out(C_s1_160));
FA FA_s1_170(.A(S_s2_170), .B(C_s2_160), .c_in(C_s3_160), .S(S_s1_170), .c_out(C_s1_170));
FA FA_s1_180(.A(S_s2_180), .B(C_s2_170), .c_in(C_s3_170), .S(S_s1_180), .c_out(C_s1_180));
FA FA_s1_190(.A(S_s2_190), .B(C_s2_180), .c_in(C_s3_180), .S(S_s1_190), .c_out(C_s1_190));
FA FA_s1_200(.A(S_s2_200), .B(C_s2_190), .c_in(C_s3_190), .S(S_s1_200), .c_out(C_s1_200));
FA FA_s1_210(.A(S_s2_210), .B(C_s2_200), .c_in(C_s3_200), .S(S_s1_210), .c_out(C_s1_210));
FA FA_s1_220(.A(S_s2_220), .B(C_s2_210), .c_in(C_s3_210), .S(S_s1_220), .c_out(C_s1_220));
FA FA_s1_230(.A(S_s2_230), .B(C_s2_220), .c_in(C_s3_220), .S(S_s1_230), .c_out(C_s1_230));
FA FA_s1_240(.A(S_s2_240), .B(C_s2_230), .c_in(C_s3_230), .S(S_s1_240), .c_out(C_s1_240));
FA FA_s1_250(.A(S_s2_250), .B(C_s2_240), .c_in(C_s3_240), .S(S_s1_250), .c_out(C_s1_250));
FA FA_s1_260(.A(S_s2_260), .B(C_s2_250), .c_in(C_s3_250), .S(S_s1_260), .c_out(C_s1_260));
FA FA_s1_270(.A(S_s2_270), .B(C_s2_260), .c_in(C_s3_260), .S(S_s1_270), .c_out(C_s1_270));
FA FA_s1_280(.A(S_s2_280), .B(C_s2_270), .c_in(C_s3_270), .S(S_s1_280), .c_out(C_s1_280));
FA FA_s1_290(.A(S_s2_290), .B(C_s2_280), .c_in(C_s3_280), .S(S_s1_290), .c_out(C_s1_290));
FA FA_s1_300(.A(S_s2_300), .B(C_s2_290), .c_in(C_s3_290), .S(S_s1_300), .c_out(C_s1_300));
FA FA_s1_310(.A(S_s2_310), .B(C_s2_300), .c_in(C_s3_300), .S(S_s1_310), .c_out(C_s1_310));
FA FA_s1_320(.A(S_s2_320), .B(C_s2_310), .c_in(C_s3_310), .S(S_s1_320), .c_out(C_s1_320));
FA FA_s1_330(.A(S_s2_330), .B(C_s2_320), .c_in(C_s3_320), .S(S_s1_330), .c_out(C_s1_330));
FA FA_s1_340(.A(S_s2_340), .B(C_s2_330), .c_in(C_s3_330), .S(S_s1_340), .c_out(C_s1_340));
FA FA_s1_350(.A(S_s2_350), .B(C_s2_340), .c_in(C_s3_340), .S(S_s1_350), .c_out(C_s1_350));
FA FA_s1_360(.A(S_s2_360), .B(C_s2_350), .c_in(C_s3_350), .S(S_s1_360), .c_out(C_s1_360));
FA FA_s1_370(.A(S_s2_370), .B(C_s2_360), .c_in(C_s3_360), .S(S_s1_370), .c_out(C_s1_370));
FA FA_s1_380(.A(S_s2_380), .B(C_s2_370), .c_in(C_s3_370), .S(S_s1_380), .c_out(C_s1_380));
FA FA_s1_390(.A(S_s2_390), .B(C_s2_380), .c_in(C_s3_380), .S(S_s1_390), .c_out(C_s1_390));
FA FA_s1_400(.A(S_s2_400), .B(C_s2_390), .c_in(C_s3_390), .S(S_s1_400), .c_out(C_s1_400));
FA FA_s1_410(.A(S_s2_410), .B(C_s2_400), .c_in(C_s3_400), .S(S_s1_410), .c_out(C_s1_410));
FA FA_s1_420(.A(S_s2_420), .B(C_s2_410), .c_in(C_s3_410), .S(S_s1_420), .c_out(C_s1_420));
FA FA_s1_430(.A(S_s2_430), .B(C_s2_420), .c_in(C_s3_420), .S(S_s1_430), .c_out(C_s1_430));
FA FA_s1_440(.A(S_s2_440), .B(C_s2_430), .c_in(C_s3_430), .S(S_s1_440), .c_out(C_s1_440));
FA FA_s1_450(.A(S_s2_450), .B(C_s2_440), .c_in(C_s3_440), .S(S_s1_450), .c_out(C_s1_450));
FA FA_s1_460(.A(S_s2_460), .B(C_s2_450), .c_in(C_s3_450), .S(S_s1_460), .c_out(C_s1_460));
FA FA_s1_470(.A(S_s2_470), .B(C_s2_460), .c_in(C_s3_460), .S(S_s1_470), .c_out(C_s1_470));
FA FA_s1_480(.A(S_s2_480), .B(C_s2_470), .c_in(C_s3_470), .S(S_s1_480), .c_out(C_s1_480));
FA FA_s1_490(.A(S_s2_490), .B(C_s2_480), .c_in(C_s3_480), .S(S_s1_490), .c_out(C_s1_490));
FA FA_s1_500(.A(S_s2_500), .B(C_s2_490), .c_in(C_s3_490), .S(S_s1_500), .c_out(C_s1_500));
FA FA_s1_510(.A(S_s2_510), .B(C_s2_500), .c_in(C_s3_500), .S(S_s1_510), .c_out(C_s1_510));
FA FA_s1_520(.A(S_s2_520), .B(C_s2_510), .c_in(C_s3_510), .S(S_s1_520), .c_out(C_s1_520));
FA FA_s1_530(.A(S_s2_530), .B(C_s2_520), .c_in(C_s3_520), .S(S_s1_530), .c_out(C_s1_530));
FA FA_s1_540(.A(S_s2_540), .B(C_s2_530), .c_in(C_s3_530), .S(S_s1_540), .c_out(C_s1_540));
FA FA_s1_550(.A(S_s2_550), .B(C_s2_540), .c_in(C_s3_540), .S(S_s1_550), .c_out(C_s1_550));
FA FA_s1_560(.A(S_s2_560), .B(C_s2_550), .c_in(C_s3_550), .S(S_s1_560), .c_out(C_s1_560));
FA FA_s1_570(.A(S_s2_570), .B(C_s2_560), .c_in(C_s3_560), .S(S_s1_570), .c_out(C_s1_570));
FA FA_s1_580(.A(S_s2_580), .B(C_s2_570), .c_in(C_s3_570), .S(S_s1_580), .c_out(C_s1_580));
FA FA_s1_590(.A(S_s2_590), .B(C_s2_580), .c_in(comb[31][28]), .S(S_s1_590), .c_out(C_s1_590));
FA FA_s1_600(.A(S_s2_600), .B(C_s2_590), .c_in(comb[31][29]), .S(S_s1_600), .c_out(C_s1_600));
FA FA_s1_610(.A(C_s2_600), .B(comb[30][31]), .c_in(comb[31][30]), .S(S_s1_610), .c_out(C_s1_610));
// stage 1 end ======================================================================= 

endmodule